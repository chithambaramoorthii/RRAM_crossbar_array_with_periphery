magic
tech sky130B
magscale 1 2
timestamp 1654740117
<< poly >>
rect 88326 435840 88526 435873
rect 88326 435670 88375 435840
rect 88477 435670 88526 435840
rect 88326 435637 88526 435670
<< polycont >>
rect 88375 435670 88477 435840
<< locali >>
rect 172220 687993 172620 688032
rect 95537 687809 95737 687969
rect 172220 687941 172259 687993
rect 172141 687861 172259 687941
rect 95437 687770 95837 687809
rect 95437 687448 95476 687770
rect 95798 687448 95837 687770
rect 120845 687623 121045 687812
rect 172140 687671 172259 687861
rect 172581 687671 172620 687993
rect 95437 687409 95837 687448
rect 120762 687584 121162 687623
rect 79772 437785 79972 437796
rect 79772 437607 79819 437785
rect 79925 437607 79972 437785
rect 79772 437596 79972 437607
rect 88326 435844 88526 435855
rect 88326 435666 88373 435844
rect 88479 435666 88526 435844
rect 80259 435645 80459 435656
rect 88326 435655 88526 435666
rect 80259 435467 80306 435645
rect 80412 435467 80459 435645
rect 80259 435456 80459 435467
rect 76602 431180 77002 431191
rect 76602 431002 76641 431180
rect 76963 431002 77002 431180
rect 76602 430991 77002 431002
rect 77400 430118 77800 430129
rect 77400 429940 77439 430118
rect 77761 429940 77800 430118
rect 77400 429929 77800 429940
rect 78409 428804 78809 428815
rect 78409 428626 78448 428804
rect 78770 428626 78809 428804
rect 78409 428615 78809 428626
rect 79436 427357 79836 427368
rect 79436 427179 79475 427357
rect 79797 427179 79836 427357
rect 79436 427168 79836 427179
rect 76601 417837 77001 417848
rect 76601 417659 76640 417837
rect 76962 417659 77001 417837
rect 76601 417648 77001 417659
rect 77400 416772 77800 416783
rect 77400 416594 77439 416772
rect 77761 416594 77800 416772
rect 77400 416583 77800 416594
rect 78411 415452 78811 415463
rect 78411 415274 78450 415452
rect 78772 415274 78811 415452
rect 78411 415263 78811 415274
rect 79435 414008 79835 414019
rect 79435 413830 79474 414008
rect 79796 413830 79835 414008
rect 79435 413819 79835 413830
rect 76602 404492 77002 404503
rect 76602 404314 76641 404492
rect 76963 404314 77002 404492
rect 76602 404303 77002 404314
rect 77400 403428 77800 403439
rect 77400 403250 77439 403428
rect 77761 403250 77800 403428
rect 77400 403239 77800 403250
rect 78409 402116 78809 402127
rect 78409 401938 78448 402116
rect 78770 401938 78809 402116
rect 78409 401927 78809 401938
rect 79435 400669 79835 400680
rect 79435 400491 79474 400669
rect 79796 400491 79835 400669
rect 79435 400480 79835 400491
rect 76602 391147 77002 391158
rect 76602 390969 76641 391147
rect 76963 390969 77002 391147
rect 76602 390958 77002 390969
rect 77400 390081 77800 390092
rect 77400 389903 77439 390081
rect 77761 389903 77800 390081
rect 77400 389892 77800 389903
rect 78409 388776 78809 388787
rect 78409 388598 78448 388776
rect 78770 388598 78809 388776
rect 78409 388587 78809 388598
rect 79430 387320 79830 387331
rect 79430 387142 79469 387320
rect 79791 387142 79830 387320
rect 79430 387131 79830 387142
rect 76602 377801 77002 377812
rect 76602 377623 76641 377801
rect 76963 377623 77002 377801
rect 76602 377612 77002 377623
rect 77400 376737 77800 376748
rect 77400 376559 77439 376737
rect 77761 376559 77800 376737
rect 77400 376548 77800 376559
rect 78409 375428 78809 375439
rect 78409 375250 78448 375428
rect 78770 375250 78809 375428
rect 78409 375239 78809 375250
rect 79434 373973 79834 373984
rect 79434 373795 79473 373973
rect 79795 373795 79834 373973
rect 79434 373784 79834 373795
rect 76601 364454 77001 364465
rect 76601 364276 76640 364454
rect 76962 364276 77001 364454
rect 76601 364265 77001 364276
rect 77400 363395 77800 363406
rect 77400 363217 77439 363395
rect 77761 363217 77800 363395
rect 77400 363206 77800 363217
rect 78406 362082 78806 362093
rect 78406 361904 78445 362082
rect 78767 361904 78806 362082
rect 78406 361893 78806 361904
rect 79436 360635 79836 360646
rect 79436 360457 79475 360635
rect 79797 360457 79836 360635
rect 79436 360446 79836 360457
rect 76601 351109 77001 351120
rect 76601 350931 76640 351109
rect 76962 350931 77001 351109
rect 76601 350920 77001 350931
rect 77400 350049 77800 350060
rect 77400 349871 77439 350049
rect 77761 349871 77800 350049
rect 77400 349860 77800 349871
rect 78409 348735 78809 348746
rect 78409 348557 78448 348735
rect 78770 348557 78809 348735
rect 78409 348546 78809 348557
rect 79435 347286 79835 347297
rect 79435 347108 79474 347286
rect 79796 347108 79835 347286
rect 79435 347097 79835 347108
rect 76601 337769 77001 337780
rect 76601 337591 76640 337769
rect 76962 337591 77001 337769
rect 76601 337580 77001 337591
rect 77400 336702 77800 336713
rect 77400 336524 77439 336702
rect 77761 336524 77800 336702
rect 77400 336513 77800 336524
rect 78404 335392 78804 335403
rect 78404 335214 78443 335392
rect 78765 335214 78804 335392
rect 78404 335203 78804 335214
rect 79435 333943 79835 333954
rect 79435 333765 79474 333943
rect 79796 333765 79835 333943
rect 79435 333754 79835 333765
rect 76602 324422 77002 324433
rect 76602 324244 76641 324422
rect 76963 324244 77002 324422
rect 76602 324233 77002 324244
rect 77400 323358 77800 323369
rect 77400 323180 77439 323358
rect 77761 323180 77800 323358
rect 77400 323169 77800 323180
rect 78409 322047 78809 322058
rect 78409 321869 78448 322047
rect 78770 321869 78809 322047
rect 78409 321858 78809 321869
rect 79438 320595 79838 320606
rect 79438 320417 79477 320595
rect 79799 320417 79838 320595
rect 79438 320406 79838 320417
rect 76600 311078 77000 311089
rect 76600 310900 76639 311078
rect 76961 310900 77000 311078
rect 76600 310889 77000 310900
rect 77400 310013 77800 310024
rect 77400 309835 77439 310013
rect 77761 309835 77800 310013
rect 77400 309824 77800 309835
rect 78410 308702 78810 308713
rect 78410 308524 78449 308702
rect 78771 308524 78810 308702
rect 78410 308513 78810 308524
rect 79431 307250 79831 307261
rect 79431 307072 79470 307250
rect 79792 307072 79831 307250
rect 79431 307061 79831 307072
rect 76602 297731 77002 297742
rect 76602 297553 76641 297731
rect 76963 297553 77002 297731
rect 76602 297542 77002 297553
rect 77400 296665 77800 296676
rect 77400 296487 77439 296665
rect 77761 296487 77800 296665
rect 77400 296476 77800 296487
rect 78411 295357 78811 295368
rect 78411 295179 78450 295357
rect 78772 295179 78811 295357
rect 78411 295168 78811 295179
rect 79437 293905 79837 293916
rect 79437 293727 79476 293905
rect 79798 293727 79837 293905
rect 79437 293716 79837 293727
rect 76602 284385 77002 284396
rect 76602 284207 76641 284385
rect 76963 284207 77002 284385
rect 76602 284196 77002 284207
rect 77400 283323 77800 283334
rect 77400 283145 77439 283323
rect 77761 283145 77800 283323
rect 77400 283134 77800 283145
rect 78409 282012 78809 282023
rect 78409 281834 78448 282012
rect 78770 281834 78809 282012
rect 78409 281823 78809 281834
rect 79433 280567 79833 280578
rect 79433 280389 79472 280567
rect 79794 280389 79833 280567
rect 79433 280378 79833 280389
rect 76601 271041 77001 271052
rect 76601 270863 76640 271041
rect 76962 270863 77001 271041
rect 76601 270852 77001 270863
rect 77400 269976 77800 269987
rect 77400 269798 77439 269976
rect 77761 269798 77800 269976
rect 77400 269787 77800 269798
rect 78410 268672 78810 268683
rect 78410 268494 78449 268672
rect 78771 268494 78810 268672
rect 78410 268483 78810 268494
rect 79436 267214 79836 267225
rect 79436 267036 79475 267214
rect 79797 267036 79836 267214
rect 79436 267025 79836 267036
rect 76601 257697 77001 257708
rect 76601 257519 76640 257697
rect 76962 257519 77001 257697
rect 76601 257508 77001 257519
rect 77400 256633 77800 256644
rect 77400 256455 77439 256633
rect 77761 256455 77800 256633
rect 77400 256444 77800 256455
rect 78409 255322 78809 255333
rect 78409 255144 78448 255322
rect 78770 255144 78809 255322
rect 78409 255133 78809 255144
rect 79436 253875 79836 253886
rect 79436 253697 79475 253875
rect 79797 253697 79836 253875
rect 79436 253686 79836 253697
rect 76602 244351 77002 244362
rect 76602 244173 76641 244351
rect 76963 244173 77002 244351
rect 76602 244162 77002 244173
rect 77400 243288 77800 243299
rect 77400 243110 77439 243288
rect 77761 243110 77800 243288
rect 77400 243099 77800 243110
rect 78411 241972 78811 241983
rect 78411 241794 78450 241972
rect 78772 241794 78811 241972
rect 78411 241783 78811 241794
rect 79437 240527 79837 240538
rect 79437 240349 79476 240527
rect 79798 240349 79837 240527
rect 79437 240338 79837 240349
rect 95537 235993 95737 687409
rect 120762 687262 120801 687584
rect 121123 687262 121162 687584
rect 146494 687501 146694 687663
rect 172140 687632 172620 687671
rect 120762 687223 121162 687262
rect 146419 687462 146819 687501
rect 120845 235980 121045 687223
rect 146419 687140 146458 687462
rect 146780 687140 146819 687462
rect 146419 687101 146819 687140
rect 146494 235981 146694 687101
rect 172140 236808 172340 687632
rect 216459 687592 216659 687845
rect 223436 687667 223636 687860
rect 223339 687628 223739 687667
rect 216358 687553 216758 687592
rect 216358 687231 216397 687553
rect 216719 687231 216758 687553
rect 223339 687306 223378 687628
rect 223700 687306 223739 687628
rect 249096 687570 249296 687811
rect 274746 687586 274946 687808
rect 300394 687622 300594 687786
rect 223339 687267 223739 687306
rect 249009 687531 249409 687570
rect 216358 687192 216758 687231
rect 203796 540602 208184 540614
rect 203796 540424 207957 540602
rect 208063 540424 208184 540602
rect 203796 540414 208184 540424
rect 207910 540413 208110 540414
rect 216459 536080 216659 687192
rect 197796 535880 216659 536080
rect 197796 235980 197996 535880
rect 223436 236473 223636 687267
rect 249009 687209 249048 687531
rect 249370 687209 249409 687531
rect 249009 687170 249409 687209
rect 274678 687547 275078 687586
rect 274678 687225 274717 687547
rect 275039 687225 275078 687547
rect 274678 687186 275078 687225
rect 300303 687583 300703 687622
rect 326043 687587 326243 687824
rect 300303 687261 300342 687583
rect 300664 687261 300703 687583
rect 300303 687222 300703 687261
rect 325939 687548 326339 687587
rect 351698 687569 351898 687902
rect 325939 687226 325978 687548
rect 326300 687226 326339 687548
rect 249096 235980 249296 687170
rect 274746 236550 274946 687186
rect 300394 236613 300594 687222
rect 325939 687187 326339 687226
rect 351604 687530 352004 687569
rect 377344 687531 377544 687736
rect 412534 687648 412734 688079
rect 412441 687609 412841 687648
rect 428648 687638 428848 687771
rect 454293 687707 454493 688308
rect 479943 687713 480143 688057
rect 454201 687668 454601 687707
rect 351604 687208 351643 687530
rect 351965 687208 352004 687530
rect 326043 236286 326243 687187
rect 351604 687169 352004 687208
rect 377265 687492 377665 687531
rect 377265 687170 377304 687492
rect 377626 687170 377665 687492
rect 412441 687287 412480 687609
rect 412802 687287 412841 687609
rect 412441 687248 412841 687287
rect 428567 687599 428967 687638
rect 428567 687277 428606 687599
rect 428928 687277 428967 687599
rect 454201 687346 454240 687668
rect 454562 687346 454601 687668
rect 454201 687307 454601 687346
rect 479850 687674 480250 687713
rect 479850 687352 479889 687674
rect 480211 687352 480250 687674
rect 479850 687313 480250 687352
rect 351698 236437 351898 687169
rect 377265 687131 377665 687170
rect 377344 235978 377544 687131
rect 412534 538574 412734 687248
rect 428567 687238 428967 687277
rect 402996 538374 412734 538574
rect 402996 235980 403196 538374
rect 428648 236395 428848 687238
rect 454293 235975 454493 687307
rect 479943 235969 480143 687313
rect 76603 230968 77003 230979
rect 76603 230790 76642 230968
rect 76964 230790 77003 230968
rect 76603 230779 77003 230790
rect 77400 229909 77800 229920
rect 77400 229731 77439 229909
rect 77761 229731 77800 229909
rect 77400 229720 77800 229731
rect 78407 228598 78807 228609
rect 78407 228420 78446 228598
rect 78768 228420 78807 228598
rect 78407 228409 78807 228420
rect 79431 227146 79831 227157
rect 79431 226968 79470 227146
rect 79792 226968 79831 227146
rect 79431 226957 79831 226968
rect 93791 216514 93991 216553
rect 93791 216192 93838 216514
rect 93944 216192 93991 216514
rect 93791 216153 93991 216192
rect 106141 216513 106341 216552
rect 106141 216191 106188 216513
rect 106294 216191 106341 216513
rect 106141 216152 106341 216191
rect 119102 216515 119302 216554
rect 119102 216193 119149 216515
rect 119255 216193 119302 216515
rect 119102 216154 119302 216193
rect 131446 216513 131646 216552
rect 131446 216191 131493 216513
rect 131599 216191 131646 216513
rect 131446 216152 131646 216191
rect 144753 216512 144953 216551
rect 144753 216190 144800 216512
rect 144906 216190 144953 216512
rect 144753 216151 144953 216190
rect 157096 216513 157296 216552
rect 157096 216191 157143 216513
rect 157249 216191 157296 216513
rect 157096 216152 157296 216191
rect 170398 216513 170598 216552
rect 170398 216191 170445 216513
rect 170551 216191 170598 216513
rect 170398 216152 170598 216191
rect 182745 216514 182945 216553
rect 182745 216192 182792 216514
rect 182898 216192 182945 216514
rect 182745 216153 182945 216192
rect 196053 216515 196253 216554
rect 196053 216193 196100 216515
rect 196206 216193 196253 216515
rect 196053 216154 196253 216193
rect 208397 216516 208597 216555
rect 208397 216194 208444 216516
rect 208550 216194 208597 216516
rect 208397 216155 208597 216194
rect 221701 216518 221901 216557
rect 221701 216196 221748 216518
rect 221854 216196 221901 216518
rect 221701 216157 221901 216196
rect 234052 216516 234252 216555
rect 234052 216194 234099 216516
rect 234205 216194 234252 216516
rect 234052 216155 234252 216194
rect 247353 216515 247553 216554
rect 247353 216193 247400 216515
rect 247506 216193 247553 216515
rect 247353 216154 247553 216193
rect 259702 216516 259902 216555
rect 259702 216194 259749 216516
rect 259855 216194 259902 216516
rect 259702 216155 259902 216194
rect 273001 216509 273201 216548
rect 273001 216187 273048 216509
rect 273154 216187 273201 216509
rect 273001 216148 273201 216187
rect 285347 216514 285547 216553
rect 285347 216192 285394 216514
rect 285500 216192 285547 216514
rect 285347 216153 285547 216192
rect 298650 216516 298850 216555
rect 298650 216194 298697 216516
rect 298803 216194 298850 216516
rect 298650 216155 298850 216194
rect 310997 216518 311197 216557
rect 310997 216196 311044 216518
rect 311150 216196 311197 216518
rect 310997 216157 311197 216196
rect 324302 216509 324502 216548
rect 324302 216187 324349 216509
rect 324455 216187 324502 216509
rect 324302 216148 324502 216187
rect 336647 216515 336847 216554
rect 336647 216193 336694 216515
rect 336800 216193 336847 216515
rect 336647 216154 336847 216193
rect 349953 216513 350153 216552
rect 349953 216191 350000 216513
rect 350106 216191 350153 216513
rect 349953 216152 350153 216191
rect 362298 216517 362498 216556
rect 362298 216195 362345 216517
rect 362451 216195 362498 216517
rect 362298 216156 362498 216195
rect 375596 216509 375796 216548
rect 375596 216187 375643 216509
rect 375749 216187 375796 216509
rect 375596 216148 375796 216187
rect 387945 216509 388145 216548
rect 387945 216187 387992 216509
rect 388098 216187 388145 216509
rect 387945 216148 388145 216187
rect 401252 216512 401452 216551
rect 401252 216190 401299 216512
rect 401405 216190 401452 216512
rect 401252 216151 401452 216190
rect 413602 216513 413802 216552
rect 413602 216191 413649 216513
rect 413755 216191 413802 216513
rect 413602 216152 413802 216191
rect 426902 216514 427102 216553
rect 426902 216192 426949 216514
rect 427055 216192 427102 216514
rect 426902 216153 427102 216192
rect 439246 216515 439446 216554
rect 439246 216193 439293 216515
rect 439399 216193 439446 216515
rect 439246 216154 439446 216193
rect 452556 216524 452756 216563
rect 452556 216202 452603 216524
rect 452709 216202 452756 216524
rect 452556 216163 452756 216202
rect 464896 216514 465096 216553
rect 464896 216192 464943 216514
rect 465049 216192 465096 216514
rect 464896 216153 465096 216192
rect 478201 216516 478401 216555
rect 478201 216194 478248 216516
rect 478354 216194 478401 216516
rect 478201 216155 478401 216194
rect 490543 216510 490743 216549
rect 490543 216188 490590 216510
rect 490696 216188 490743 216510
rect 490543 216149 490743 216188
rect 94848 215760 95048 215799
rect 94848 215438 94895 215760
rect 95001 215438 95048 215760
rect 94848 215399 95048 215438
rect 107198 215760 107398 215799
rect 107198 215438 107245 215760
rect 107351 215438 107398 215760
rect 107198 215399 107398 215438
rect 120163 215760 120363 215799
rect 120163 215438 120210 215760
rect 120316 215438 120363 215760
rect 120163 215399 120363 215438
rect 132507 215757 132707 215796
rect 132507 215435 132554 215757
rect 132660 215435 132707 215757
rect 132507 215396 132707 215435
rect 145814 215760 146014 215799
rect 145814 215438 145861 215760
rect 145967 215438 146014 215760
rect 145814 215399 146014 215438
rect 158154 215753 158354 215792
rect 158154 215431 158201 215753
rect 158307 215431 158354 215753
rect 158154 215392 158354 215431
rect 171464 215759 171664 215798
rect 171464 215437 171511 215759
rect 171617 215437 171664 215759
rect 171464 215398 171664 215437
rect 183807 215760 184007 215799
rect 183807 215438 183854 215760
rect 183960 215438 184007 215760
rect 183807 215399 184007 215438
rect 197110 215761 197310 215800
rect 197110 215439 197157 215761
rect 197263 215439 197310 215761
rect 197110 215400 197310 215439
rect 209458 215761 209658 215800
rect 209458 215439 209505 215761
rect 209611 215439 209658 215761
rect 209458 215400 209658 215439
rect 222764 215761 222964 215800
rect 222764 215439 222811 215761
rect 222917 215439 222964 215761
rect 222764 215400 222964 215439
rect 235107 215761 235307 215800
rect 235107 215439 235154 215761
rect 235260 215439 235307 215761
rect 235107 215400 235307 215439
rect 248409 215760 248609 215799
rect 248409 215438 248456 215760
rect 248562 215438 248609 215760
rect 248409 215399 248609 215438
rect 260760 215761 260960 215800
rect 260760 215439 260807 215761
rect 260913 215439 260960 215761
rect 260760 215400 260960 215439
rect 274061 215759 274261 215798
rect 274061 215437 274108 215759
rect 274214 215437 274261 215759
rect 274061 215398 274261 215437
rect 286405 215759 286605 215798
rect 286405 215437 286452 215759
rect 286558 215437 286605 215759
rect 286405 215398 286605 215437
rect 299709 215761 299909 215800
rect 299709 215439 299756 215761
rect 299862 215439 299909 215761
rect 299709 215400 299909 215439
rect 312056 215761 312256 215800
rect 312056 215439 312103 215761
rect 312209 215439 312256 215761
rect 312056 215400 312256 215439
rect 325361 215759 325561 215798
rect 325361 215437 325408 215759
rect 325514 215437 325561 215759
rect 325361 215398 325561 215437
rect 337706 215756 337906 215795
rect 337706 215434 337753 215756
rect 337859 215434 337906 215756
rect 337706 215395 337906 215434
rect 351008 215759 351208 215798
rect 351008 215437 351055 215759
rect 351161 215437 351208 215759
rect 351008 215398 351208 215437
rect 363357 215759 363557 215798
rect 363357 215437 363404 215759
rect 363510 215437 363557 215759
rect 363357 215398 363557 215437
rect 376662 215756 376862 215795
rect 376662 215434 376709 215756
rect 376815 215434 376862 215756
rect 376662 215395 376862 215434
rect 389004 215762 389204 215801
rect 389004 215440 389051 215762
rect 389157 215440 389204 215762
rect 389004 215401 389204 215440
rect 402311 215758 402511 215797
rect 402311 215436 402358 215758
rect 402464 215436 402511 215758
rect 402311 215397 402511 215436
rect 414658 215756 414858 215795
rect 414658 215434 414705 215756
rect 414811 215434 414858 215756
rect 414658 215395 414858 215434
rect 427961 215763 428161 215802
rect 427961 215441 428008 215763
rect 428114 215441 428161 215763
rect 427961 215402 428161 215441
rect 440306 215757 440506 215796
rect 440306 215435 440353 215757
rect 440459 215435 440506 215757
rect 440306 215396 440506 215435
rect 453612 215763 453812 215802
rect 453612 215441 453659 215763
rect 453765 215441 453812 215763
rect 453612 215402 453812 215441
rect 465958 215761 466158 215800
rect 465958 215439 466005 215761
rect 466111 215439 466158 215761
rect 465958 215400 466158 215439
rect 479259 215759 479459 215798
rect 479259 215437 479306 215759
rect 479412 215437 479459 215759
rect 479259 215398 479459 215437
rect 491606 215759 491806 215798
rect 491606 215437 491653 215759
rect 491759 215437 491806 215759
rect 491606 215398 491806 215437
rect 96165 214879 96365 214918
rect 96165 214557 96212 214879
rect 96318 214557 96365 214879
rect 96165 214518 96365 214557
rect 108508 214882 108708 214921
rect 108508 214560 108555 214882
rect 108661 214560 108708 214882
rect 108508 214521 108708 214560
rect 121474 214876 121674 214915
rect 121474 214554 121521 214876
rect 121627 214554 121674 214876
rect 121474 214515 121674 214554
rect 133818 214878 134018 214917
rect 133818 214556 133865 214878
rect 133971 214556 134018 214878
rect 133818 214517 134018 214556
rect 147122 214878 147322 214917
rect 147122 214556 147169 214878
rect 147275 214556 147322 214878
rect 147122 214517 147322 214556
rect 159470 214881 159670 214920
rect 159470 214559 159517 214881
rect 159623 214559 159670 214881
rect 159470 214520 159670 214559
rect 172774 214879 172974 214918
rect 172774 214557 172821 214879
rect 172927 214557 172974 214879
rect 172774 214518 172974 214557
rect 185121 214879 185321 214918
rect 185121 214557 185168 214879
rect 185274 214557 185321 214879
rect 185121 214518 185321 214557
rect 198422 214877 198622 214916
rect 198422 214555 198469 214877
rect 198575 214555 198622 214877
rect 198422 214516 198622 214555
rect 210771 214878 210971 214917
rect 210771 214556 210818 214878
rect 210924 214556 210971 214878
rect 210771 214517 210971 214556
rect 224078 214881 224278 214920
rect 224078 214559 224125 214881
rect 224231 214559 224278 214881
rect 224078 214520 224278 214559
rect 236418 214879 236618 214918
rect 236418 214557 236465 214879
rect 236571 214557 236618 214879
rect 236418 214518 236618 214557
rect 249722 214876 249922 214915
rect 249722 214554 249769 214876
rect 249875 214554 249922 214876
rect 249722 214515 249922 214554
rect 262070 214880 262270 214919
rect 262070 214558 262117 214880
rect 262223 214558 262270 214880
rect 262070 214519 262270 214558
rect 275373 214878 275573 214917
rect 275373 214556 275420 214878
rect 275526 214556 275573 214878
rect 275373 214517 275573 214556
rect 287721 214878 287921 214917
rect 287721 214556 287768 214878
rect 287874 214556 287921 214878
rect 287721 214517 287921 214556
rect 301030 214881 301230 214920
rect 301030 214559 301077 214881
rect 301183 214559 301230 214881
rect 301030 214520 301230 214559
rect 313368 214879 313568 214918
rect 313368 214557 313415 214879
rect 313521 214557 313568 214879
rect 313368 214518 313568 214557
rect 326673 214878 326873 214917
rect 326673 214556 326720 214878
rect 326826 214556 326873 214878
rect 326673 214517 326873 214556
rect 339018 214879 339218 214918
rect 339018 214557 339065 214879
rect 339171 214557 339218 214879
rect 339018 214518 339218 214557
rect 352324 214876 352524 214915
rect 352324 214554 352371 214876
rect 352477 214554 352524 214876
rect 352324 214515 352524 214554
rect 364669 214879 364869 214918
rect 364669 214557 364716 214879
rect 364822 214557 364869 214879
rect 364669 214518 364869 214557
rect 377974 214879 378174 214918
rect 377974 214557 378021 214879
rect 378127 214557 378174 214879
rect 377974 214518 378174 214557
rect 390321 214877 390521 214916
rect 390321 214555 390368 214877
rect 390474 214555 390521 214877
rect 390321 214516 390521 214555
rect 403614 214869 403814 214908
rect 403614 214547 403661 214869
rect 403767 214547 403814 214869
rect 403614 214508 403814 214547
rect 415966 214873 416166 214912
rect 415966 214551 416013 214873
rect 416119 214551 416166 214873
rect 415966 214512 416166 214551
rect 429276 214876 429476 214915
rect 429276 214554 429323 214876
rect 429429 214554 429476 214876
rect 429276 214515 429476 214554
rect 441618 214879 441818 214918
rect 441618 214557 441665 214879
rect 441771 214557 441818 214879
rect 441618 214518 441818 214557
rect 454924 214882 455124 214921
rect 454924 214560 454971 214882
rect 455077 214560 455124 214882
rect 454924 214521 455124 214560
rect 467268 214877 467468 214916
rect 467268 214555 467315 214877
rect 467421 214555 467468 214877
rect 467268 214516 467468 214555
rect 480569 214876 480769 214915
rect 480569 214554 480616 214876
rect 480722 214554 480769 214876
rect 480569 214515 480769 214554
rect 492922 214877 493122 214916
rect 492922 214555 492969 214877
rect 493075 214555 493122 214877
rect 492922 214516 493122 214555
rect 97613 214090 97813 214129
rect 97613 213768 97660 214090
rect 97766 213768 97813 214090
rect 97613 213729 97813 213768
rect 109971 214086 110171 214125
rect 109971 213764 110018 214086
rect 110124 213764 110171 214086
rect 109971 213725 110171 213764
rect 122925 214091 123125 214130
rect 122925 213769 122972 214091
rect 123078 213769 123125 214091
rect 122925 213730 123125 213769
rect 135288 214088 135488 214127
rect 135288 213766 135335 214088
rect 135441 213766 135488 214088
rect 135288 213727 135488 213766
rect 148581 214080 148781 214119
rect 148581 213758 148628 214080
rect 148734 213758 148781 214080
rect 148581 213719 148781 213758
rect 160921 214080 161121 214119
rect 160921 213758 160968 214080
rect 161074 213758 161121 214080
rect 160921 213719 161121 213758
rect 174225 214086 174425 214125
rect 174225 213764 174272 214086
rect 174378 213764 174425 214086
rect 174225 213725 174425 213764
rect 186585 214098 186785 214137
rect 186585 213776 186632 214098
rect 186738 213776 186785 214098
rect 186585 213737 186785 213776
rect 199877 214080 200077 214119
rect 199877 213758 199924 214080
rect 200030 213758 200077 214080
rect 199877 213719 200077 213758
rect 212226 214094 212426 214133
rect 212226 213772 212273 214094
rect 212379 213772 212426 214094
rect 212226 213733 212426 213772
rect 225532 214088 225732 214127
rect 225532 213766 225579 214088
rect 225685 213766 225732 214088
rect 225532 213727 225732 213766
rect 237886 214090 238086 214129
rect 237886 213768 237933 214090
rect 238039 213768 238086 214090
rect 237886 213729 238086 213768
rect 251189 214091 251389 214130
rect 251189 213769 251236 214091
rect 251342 213769 251389 214091
rect 251189 213730 251389 213769
rect 263531 214095 263731 214134
rect 263531 213773 263578 214095
rect 263684 213773 263731 214095
rect 263531 213734 263731 213773
rect 276838 214086 277038 214125
rect 276838 213764 276885 214086
rect 276991 213764 277038 214086
rect 276838 213725 277038 213764
rect 289167 214085 289367 214124
rect 289167 213763 289214 214085
rect 289320 213763 289367 214085
rect 289167 213724 289367 213763
rect 302486 214088 302686 214127
rect 302486 213766 302533 214088
rect 302639 213766 302686 214088
rect 302486 213727 302686 213766
rect 314825 214091 315025 214130
rect 314825 213769 314872 214091
rect 314978 213769 315025 214091
rect 314825 213730 315025 213769
rect 328123 214091 328323 214130
rect 328123 213769 328170 214091
rect 328276 213769 328323 214091
rect 328123 213730 328323 213769
rect 340473 214092 340673 214131
rect 340473 213770 340520 214092
rect 340626 213770 340673 214092
rect 340473 213731 340673 213770
rect 353782 214088 353982 214127
rect 353782 213766 353829 214088
rect 353935 213766 353982 214088
rect 353782 213727 353982 213766
rect 366116 214093 366316 214132
rect 366116 213771 366163 214093
rect 366269 213771 366316 214093
rect 366116 213732 366316 213771
rect 379434 214092 379634 214131
rect 379434 213770 379481 214092
rect 379587 213770 379634 214092
rect 379434 213731 379634 213770
rect 391768 214089 391968 214128
rect 391768 213767 391815 214089
rect 391921 213767 391968 214089
rect 391768 213728 391968 213767
rect 405079 214085 405279 214124
rect 405079 213763 405126 214085
rect 405232 213763 405279 214085
rect 405079 213724 405279 213763
rect 417427 214095 417627 214134
rect 417427 213773 417474 214095
rect 417580 213773 417627 214095
rect 417427 213734 417627 213773
rect 430742 214094 430942 214133
rect 430742 213772 430789 214094
rect 430895 213772 430942 214094
rect 430742 213733 430942 213772
rect 443078 214088 443278 214127
rect 443078 213766 443125 214088
rect 443231 213766 443278 214088
rect 443078 213727 443278 213766
rect 456383 214088 456583 214127
rect 456383 213766 456430 214088
rect 456536 213766 456583 214088
rect 456383 213727 456583 213766
rect 468736 214094 468936 214133
rect 468736 213772 468783 214094
rect 468889 213772 468936 214094
rect 468736 213733 468936 213772
rect 482038 214088 482238 214127
rect 482038 213766 482085 214088
rect 482191 213766 482238 214088
rect 482038 213727 482238 213766
rect 494373 214089 494573 214128
rect 494373 213767 494420 214089
rect 494526 213767 494573 214089
rect 494373 213728 494573 213767
<< viali >>
rect 95476 687448 95798 687770
rect 172259 687671 172581 687993
rect 79819 437607 79925 437785
rect 88373 435840 88479 435844
rect 88373 435670 88375 435840
rect 88375 435670 88477 435840
rect 88477 435670 88479 435840
rect 88373 435666 88479 435670
rect 80306 435467 80412 435645
rect 76641 431002 76963 431180
rect 77439 429940 77761 430118
rect 78448 428626 78770 428804
rect 79475 427179 79797 427357
rect 76640 417659 76962 417837
rect 77439 416594 77761 416772
rect 78450 415274 78772 415452
rect 79474 413830 79796 414008
rect 76641 404314 76963 404492
rect 77439 403250 77761 403428
rect 78448 401938 78770 402116
rect 79474 400491 79796 400669
rect 76641 390969 76963 391147
rect 77439 389903 77761 390081
rect 78448 388598 78770 388776
rect 79469 387142 79791 387320
rect 76641 377623 76963 377801
rect 77439 376559 77761 376737
rect 78448 375250 78770 375428
rect 79473 373795 79795 373973
rect 76640 364276 76962 364454
rect 77439 363217 77761 363395
rect 78445 361904 78767 362082
rect 79475 360457 79797 360635
rect 76640 350931 76962 351109
rect 77439 349871 77761 350049
rect 78448 348557 78770 348735
rect 79474 347108 79796 347286
rect 76640 337591 76962 337769
rect 77439 336524 77761 336702
rect 78443 335214 78765 335392
rect 79474 333765 79796 333943
rect 76641 324244 76963 324422
rect 77439 323180 77761 323358
rect 78448 321869 78770 322047
rect 79477 320417 79799 320595
rect 76639 310900 76961 311078
rect 77439 309835 77761 310013
rect 78449 308524 78771 308702
rect 79470 307072 79792 307250
rect 76641 297553 76963 297731
rect 77439 296487 77761 296665
rect 78450 295179 78772 295357
rect 79476 293727 79798 293905
rect 76641 284207 76963 284385
rect 77439 283145 77761 283323
rect 78448 281834 78770 282012
rect 79472 280389 79794 280567
rect 76640 270863 76962 271041
rect 77439 269798 77761 269976
rect 78449 268494 78771 268672
rect 79475 267036 79797 267214
rect 76640 257519 76962 257697
rect 77439 256455 77761 256633
rect 78448 255144 78770 255322
rect 79475 253697 79797 253875
rect 76641 244173 76963 244351
rect 77439 243110 77761 243288
rect 78450 241794 78772 241972
rect 79476 240349 79798 240527
rect 120801 687262 121123 687584
rect 146458 687140 146780 687462
rect 216397 687231 216719 687553
rect 223378 687306 223700 687628
rect 207957 540424 208063 540602
rect 249048 687209 249370 687531
rect 274717 687225 275039 687547
rect 300342 687261 300664 687583
rect 325978 687226 326300 687548
rect 351643 687208 351965 687530
rect 377304 687170 377626 687492
rect 412480 687287 412802 687609
rect 428606 687277 428928 687599
rect 454240 687346 454562 687668
rect 479889 687352 480211 687674
rect 76642 230790 76964 230968
rect 77439 229731 77761 229909
rect 78446 228420 78768 228598
rect 79470 226968 79792 227146
rect 93838 216192 93944 216514
rect 106188 216191 106294 216513
rect 119149 216193 119255 216515
rect 131493 216191 131599 216513
rect 144800 216190 144906 216512
rect 157143 216191 157249 216513
rect 170445 216191 170551 216513
rect 182792 216192 182898 216514
rect 196100 216193 196206 216515
rect 208444 216194 208550 216516
rect 221748 216196 221854 216518
rect 234099 216194 234205 216516
rect 247400 216193 247506 216515
rect 259749 216194 259855 216516
rect 273048 216187 273154 216509
rect 285394 216192 285500 216514
rect 298697 216194 298803 216516
rect 311044 216196 311150 216518
rect 324349 216187 324455 216509
rect 336694 216193 336800 216515
rect 350000 216191 350106 216513
rect 362345 216195 362451 216517
rect 375643 216187 375749 216509
rect 387992 216187 388098 216509
rect 401299 216190 401405 216512
rect 413649 216191 413755 216513
rect 426949 216192 427055 216514
rect 439293 216193 439399 216515
rect 452603 216202 452709 216524
rect 464943 216192 465049 216514
rect 478248 216194 478354 216516
rect 490590 216188 490696 216510
rect 94895 215438 95001 215760
rect 107245 215438 107351 215760
rect 120210 215438 120316 215760
rect 132554 215435 132660 215757
rect 145861 215438 145967 215760
rect 158201 215431 158307 215753
rect 171511 215437 171617 215759
rect 183854 215438 183960 215760
rect 197157 215439 197263 215761
rect 209505 215439 209611 215761
rect 222811 215439 222917 215761
rect 235154 215439 235260 215761
rect 248456 215438 248562 215760
rect 260807 215439 260913 215761
rect 274108 215437 274214 215759
rect 286452 215437 286558 215759
rect 299756 215439 299862 215761
rect 312103 215439 312209 215761
rect 325408 215437 325514 215759
rect 337753 215434 337859 215756
rect 351055 215437 351161 215759
rect 363404 215437 363510 215759
rect 376709 215434 376815 215756
rect 389051 215440 389157 215762
rect 402358 215436 402464 215758
rect 414705 215434 414811 215756
rect 428008 215441 428114 215763
rect 440353 215435 440459 215757
rect 453659 215441 453765 215763
rect 466005 215439 466111 215761
rect 479306 215437 479412 215759
rect 491653 215437 491759 215759
rect 96212 214557 96318 214879
rect 108555 214560 108661 214882
rect 121521 214554 121627 214876
rect 133865 214556 133971 214878
rect 147169 214556 147275 214878
rect 159517 214559 159623 214881
rect 172821 214557 172927 214879
rect 185168 214557 185274 214879
rect 198469 214555 198575 214877
rect 210818 214556 210924 214878
rect 224125 214559 224231 214881
rect 236465 214557 236571 214879
rect 249769 214554 249875 214876
rect 262117 214558 262223 214880
rect 275420 214556 275526 214878
rect 287768 214556 287874 214878
rect 301077 214559 301183 214881
rect 313415 214557 313521 214879
rect 326720 214556 326826 214878
rect 339065 214557 339171 214879
rect 352371 214554 352477 214876
rect 364716 214557 364822 214879
rect 378021 214557 378127 214879
rect 390368 214555 390474 214877
rect 403661 214547 403767 214869
rect 416013 214551 416119 214873
rect 429323 214554 429429 214876
rect 441665 214557 441771 214879
rect 454971 214560 455077 214882
rect 467315 214555 467421 214877
rect 480616 214554 480722 214876
rect 492969 214555 493075 214877
rect 97660 213768 97766 214090
rect 110018 213764 110124 214086
rect 122972 213769 123078 214091
rect 135335 213766 135441 214088
rect 148628 213758 148734 214080
rect 160968 213758 161074 214080
rect 174272 213764 174378 214086
rect 186632 213776 186738 214098
rect 199924 213758 200030 214080
rect 212273 213772 212379 214094
rect 225579 213766 225685 214088
rect 237933 213768 238039 214090
rect 251236 213769 251342 214091
rect 263578 213773 263684 214095
rect 276885 213764 276991 214086
rect 289214 213763 289320 214085
rect 302533 213766 302639 214088
rect 314872 213769 314978 214091
rect 328170 213769 328276 214091
rect 340520 213770 340626 214092
rect 353829 213766 353935 214088
rect 366163 213771 366269 214093
rect 379481 213770 379587 214092
rect 391815 213767 391921 214089
rect 405126 213763 405232 214085
rect 417474 213773 417580 214095
rect 430789 213772 430895 214094
rect 443125 213766 443231 214088
rect 456430 213766 456536 214088
rect 468783 213772 468889 214094
rect 482085 213766 482191 214088
rect 494420 213767 494526 214089
<< metal1 >>
rect 172220 688018 172620 688032
rect 95437 687795 95837 687809
rect 95437 687423 95451 687795
rect 95823 687423 95837 687795
rect 172220 687646 172234 688018
rect 172606 687646 172620 688018
rect 454201 687693 454601 687707
rect 172220 687632 172620 687646
rect 223339 687653 223739 687667
rect 95437 687409 95837 687423
rect 120762 687609 121162 687623
rect 120762 687237 120776 687609
rect 121148 687237 121162 687609
rect 216358 687578 216758 687592
rect 120762 687223 121162 687237
rect 146419 687487 146819 687501
rect 146419 687115 146433 687487
rect 146805 687115 146819 687487
rect 216358 687206 216372 687578
rect 216744 687206 216758 687578
rect 223339 687281 223353 687653
rect 223725 687281 223739 687653
rect 412441 687634 412841 687648
rect 300303 687608 300703 687622
rect 274678 687572 275078 687586
rect 223339 687267 223739 687281
rect 249009 687556 249409 687570
rect 216358 687192 216758 687206
rect 249009 687184 249023 687556
rect 249395 687184 249409 687556
rect 274678 687200 274692 687572
rect 275064 687200 275078 687572
rect 300303 687236 300317 687608
rect 300689 687236 300703 687608
rect 300303 687222 300703 687236
rect 325939 687573 326339 687587
rect 274678 687186 275078 687200
rect 325939 687201 325953 687573
rect 326325 687201 326339 687573
rect 325939 687187 326339 687201
rect 351604 687555 352004 687569
rect 249009 687170 249409 687184
rect 351604 687183 351618 687555
rect 351990 687183 352004 687555
rect 351604 687169 352004 687183
rect 377265 687517 377665 687531
rect 377265 687145 377279 687517
rect 377651 687145 377665 687517
rect 412441 687262 412455 687634
rect 412827 687262 412841 687634
rect 412441 687248 412841 687262
rect 428567 687624 428967 687638
rect 428567 687252 428581 687624
rect 428953 687252 428967 687624
rect 454201 687321 454215 687693
rect 454587 687321 454601 687693
rect 454201 687307 454601 687321
rect 479850 687699 480250 687713
rect 479850 687327 479864 687699
rect 480236 687327 480250 687699
rect 479850 687313 480250 687327
rect 428567 687238 428967 687252
rect 377265 687131 377665 687145
rect 146419 687101 146819 687115
rect 189821 660815 190221 660853
rect 189821 660801 190222 660815
rect 189821 660429 189836 660801
rect 190208 660429 190222 660801
rect 189821 660415 190222 660429
rect 189821 549806 190221 660415
rect 207910 601904 569346 601914
rect 207910 601724 569028 601904
rect 569208 601724 569346 601904
rect 207910 601714 569346 601724
rect 204005 557076 206574 557276
rect 197183 550264 197383 550274
rect 197183 550084 197193 550264
rect 197373 550084 197383 550264
rect 197183 550074 197383 550084
rect 200939 550264 201139 550274
rect 200939 550084 200949 550264
rect 201129 550084 201139 550264
rect 200939 550074 201139 550084
rect 200934 548989 201134 548999
rect 200934 548809 200944 548989
rect 201124 548809 201134 548989
rect 200934 548799 201134 548809
rect 193931 548533 194131 548543
rect 193931 548353 193941 548533
rect 194121 548353 194131 548533
rect 193931 548343 194131 548353
rect 199418 548378 199780 548406
rect 199418 548198 199445 548378
rect 199753 548198 199780 548378
rect 199418 548170 199780 548198
rect 193007 539403 193207 540649
rect 196618 539911 196818 540728
rect 198268 539911 198468 540705
rect 196618 539901 198468 539911
rect 196618 539721 198062 539901
rect 198242 539721 198468 539901
rect 196618 539711 198468 539721
rect 201925 539403 202125 540634
rect 193007 539393 202125 539403
rect 193007 539213 201881 539393
rect 202061 539213 202125 539393
rect 193007 539203 202125 539213
rect 206374 530912 206574 557076
rect 207910 540602 208110 601714
rect 207910 540424 207957 540602
rect 208063 540424 208110 540602
rect 207910 540413 208110 540424
rect 208749 600903 565743 600913
rect 208749 600723 565481 600903
rect 565661 600723 565743 600903
rect 208749 600713 565743 600723
rect 208749 539899 208949 600713
rect 208749 539719 208759 539899
rect 208939 539719 208949 539899
rect 208749 539709 208949 539719
rect 209972 599648 562162 599659
rect 209972 599468 561939 599648
rect 562119 599468 562162 599648
rect 209972 599459 562162 599468
rect 209972 539393 210172 599459
rect 561929 599458 562129 599459
rect 417736 577766 558642 577776
rect 417736 577765 558400 577766
rect 417736 577585 417834 577765
rect 418014 577586 558400 577765
rect 558580 577586 558642 577766
rect 418014 577585 558642 577586
rect 417736 577576 558642 577585
rect 417824 577575 418024 577576
rect 417759 577176 555088 577186
rect 417759 576996 417838 577176
rect 418018 576996 554850 577176
rect 555030 576996 555088 577176
rect 417759 576986 555088 576996
rect 417754 576449 551552 576459
rect 417754 576269 417861 576449
rect 418041 576269 551301 576449
rect 551481 576269 551552 576449
rect 417754 576259 551552 576269
rect 410946 557128 422249 557328
rect 404128 550381 404328 550391
rect 396661 550225 397240 550362
rect 396661 550045 396874 550225
rect 397054 550045 397240 550225
rect 404128 550201 404138 550381
rect 404318 550201 404328 550381
rect 404128 550191 404328 550201
rect 407882 550382 408082 550392
rect 407882 550202 407892 550382
rect 408072 550202 408082 550382
rect 407882 550192 408082 550202
rect 396661 549892 397240 550045
rect 406476 548434 406728 548460
rect 406476 548254 406512 548434
rect 406692 548254 406728 548434
rect 406476 548228 406728 548254
rect 209972 539213 209982 539393
rect 210162 539213 210172 539393
rect 399962 539569 400162 540718
rect 403575 540021 403775 540791
rect 405227 540021 405427 540764
rect 403575 540011 405427 540021
rect 403575 539831 405237 540011
rect 405417 539831 405427 540011
rect 403575 539821 405427 539831
rect 408860 539569 409060 540701
rect 399962 539559 409060 539569
rect 399962 539379 408870 539559
rect 409050 539379 409060 539559
rect 399962 539369 409060 539379
rect 209972 539203 210172 539213
rect 206374 530732 206384 530912
rect 206564 530732 206574 530912
rect 206374 530722 206574 530732
rect 422049 530923 422249 557128
rect 422049 530913 422250 530923
rect 422049 530733 422060 530913
rect 422240 530733 422250 530913
rect 422049 530724 422250 530733
rect 422050 530723 422250 530724
rect 300899 525619 301099 525629
rect 300899 525439 300909 525619
rect 301089 525439 301099 525619
rect 300899 525429 301099 525439
rect 480462 520790 480662 520800
rect 480462 520610 480472 520790
rect 480652 520610 480662 520790
rect 480462 520600 480662 520610
rect 275058 519734 275572 519744
rect 275058 519234 275097 519734
rect 275533 519234 275572 519734
rect 275058 519224 275572 519234
rect 326549 518225 326749 518235
rect 326549 518045 326559 518225
rect 326739 518045 326749 518225
rect 326549 518035 326749 518045
rect 352199 510797 352399 510807
rect 352199 510617 352209 510797
rect 352389 510617 352399 510797
rect 352199 510607 352399 510617
rect 454799 510596 454999 510606
rect 454799 510416 454809 510596
rect 454989 510416 454999 510596
rect 454799 510406 454999 510416
rect 377857 503373 378057 503383
rect 377857 503193 377867 503373
rect 378047 503193 378057 503373
rect 377857 503183 378057 503193
rect 429152 503211 429352 503221
rect 429152 503031 429162 503211
rect 429342 503031 429352 503211
rect 429152 503021 429352 503031
rect 407257 494410 407457 494420
rect 407257 494230 407267 494410
rect 407447 494230 407457 494410
rect 407257 494220 407457 494230
rect 95989 446131 96189 446141
rect 95989 445951 95999 446131
rect 96179 445951 96189 446131
rect 95989 445941 96189 445951
rect 75882 437847 76063 438069
rect 76124 438045 76324 438055
rect 76124 437865 76134 438045
rect 76314 437865 76324 438045
rect 76124 437855 76324 437865
rect 79772 437786 79972 437796
rect 79772 437606 79782 437786
rect 79962 437606 79972 437786
rect 79772 437596 79972 437606
rect 40073 436045 76002 436145
rect 40073 42884 40173 436045
rect 88326 435845 88526 435855
rect 88326 435665 88336 435845
rect 88516 435665 88526 435845
rect 80259 435646 80459 435656
rect 88326 435655 88526 435665
rect 80259 435466 80269 435646
rect 80449 435466 80459 435646
rect 80259 435456 80459 435466
rect 76141 435289 76341 435299
rect 76141 435109 76151 435289
rect 76331 435109 76341 435289
rect 76141 435099 76341 435109
rect 77072 434133 77272 434143
rect 77072 433953 77082 434133
rect 77262 433953 77272 434133
rect 77072 433943 77272 433953
rect 79003 433185 79203 433195
rect 79003 433005 79013 433185
rect 79193 433005 79203 433185
rect 79003 432995 79203 433005
rect 75878 430875 76226 431345
rect 76602 431181 77002 431191
rect 76602 431001 76616 431181
rect 76988 431001 77002 431181
rect 76602 430991 77002 431001
rect 75876 429753 76270 430279
rect 77400 430119 77800 430129
rect 77400 429939 77414 430119
rect 77786 429939 77800 430119
rect 77400 429929 77800 429939
rect 75892 428471 76262 428979
rect 78409 428805 78809 428815
rect 78409 428625 78423 428805
rect 78795 428625 78809 428805
rect 78409 428615 78809 428625
rect 75890 426989 76352 427501
rect 79436 427358 79836 427368
rect 79436 427178 79450 427358
rect 79822 427178 79836 427358
rect 79436 427168 79836 427178
rect 76151 424705 76351 424715
rect 76151 424525 76161 424705
rect 76341 424525 76351 424705
rect 76151 424515 76351 424525
rect 40584 422678 76008 422778
rect 40584 43186 40684 422678
rect 76166 421939 76366 421949
rect 76166 421759 76176 421939
rect 76356 421759 76366 421939
rect 76166 421749 76366 421759
rect 77105 420781 77305 420791
rect 77105 420601 77115 420781
rect 77295 420601 77305 420781
rect 77105 420591 77305 420601
rect 78994 419838 79194 419848
rect 78994 419658 79004 419838
rect 79184 419658 79194 419838
rect 78994 419648 79194 419658
rect 76601 417838 77001 417848
rect 76601 417658 76615 417838
rect 76987 417658 77001 417838
rect 76601 417648 77001 417658
rect 77400 416773 77800 416783
rect 77400 416593 77414 416773
rect 77786 416593 77800 416773
rect 77400 416583 77800 416593
rect 78411 415453 78811 415463
rect 78411 415273 78425 415453
rect 78797 415273 78811 415453
rect 78411 415263 78811 415273
rect 79435 414009 79835 414019
rect 79435 413829 79449 414009
rect 79821 413829 79835 414009
rect 79435 413819 79835 413829
rect 76135 411361 76335 411371
rect 76135 411181 76145 411361
rect 76325 411181 76335 411361
rect 76135 411171 76335 411181
rect 41051 409345 76005 409445
rect 41051 43404 41151 409345
rect 76166 408594 76366 408604
rect 76166 408414 76176 408594
rect 76356 408414 76366 408594
rect 76166 408404 76366 408414
rect 77093 407441 77293 407451
rect 77093 407261 77103 407441
rect 77283 407261 77293 407441
rect 77093 407251 77293 407261
rect 78978 406493 79178 406503
rect 78978 406313 78988 406493
rect 79168 406313 79178 406493
rect 78978 406303 79178 406313
rect 76602 404493 77002 404503
rect 76602 404313 76616 404493
rect 76988 404313 77002 404493
rect 76602 404303 77002 404313
rect 77400 403429 77800 403439
rect 77400 403249 77414 403429
rect 77786 403249 77800 403429
rect 77400 403239 77800 403249
rect 78409 402117 78809 402127
rect 78409 401937 78423 402117
rect 78795 401937 78809 402117
rect 78409 401927 78809 401937
rect 79435 400670 79835 400680
rect 79435 400490 79449 400670
rect 79821 400490 79835 400670
rect 79435 400480 79835 400490
rect 76148 398006 76348 398016
rect 76148 397826 76158 398006
rect 76338 397826 76348 398006
rect 76148 397816 76348 397826
rect 41558 395993 75998 396093
rect 41558 47261 41658 395993
rect 76153 395252 76353 395262
rect 76153 395072 76163 395252
rect 76343 395072 76353 395252
rect 76153 395062 76353 395072
rect 77105 394092 77305 394102
rect 77105 393912 77115 394092
rect 77295 393912 77305 394092
rect 77105 393902 77305 393912
rect 79003 393153 79203 393163
rect 79003 392973 79013 393153
rect 79193 392973 79203 393153
rect 79003 392963 79203 392973
rect 76602 391148 77002 391158
rect 76602 390968 76616 391148
rect 76988 390968 77002 391148
rect 76602 390958 77002 390968
rect 77400 390082 77800 390092
rect 77400 389902 77414 390082
rect 77786 389902 77800 390082
rect 77400 389892 77800 389902
rect 78409 388777 78809 388787
rect 78409 388597 78423 388777
rect 78795 388597 78809 388777
rect 78409 388587 78809 388597
rect 79430 387321 79830 387331
rect 79430 387141 79444 387321
rect 79816 387141 79830 387321
rect 79430 387131 79830 387141
rect 76123 384666 76323 384676
rect 76123 384486 76133 384666
rect 76313 384486 76323 384666
rect 76123 384476 76323 384486
rect 42172 382649 75996 382749
rect 41558 47257 41659 47261
rect 41559 43646 41659 47257
rect 42172 43878 42272 382649
rect 76128 381904 76328 381914
rect 76128 381724 76138 381904
rect 76318 381724 76328 381904
rect 76128 381714 76328 381724
rect 77093 380748 77293 380758
rect 77093 380568 77103 380748
rect 77283 380568 77293 380748
rect 77093 380558 77293 380568
rect 78969 379806 79169 379816
rect 78969 379626 78979 379806
rect 79159 379626 79169 379806
rect 78969 379616 79169 379626
rect 76602 377802 77002 377812
rect 76602 377622 76616 377802
rect 76988 377622 77002 377802
rect 76602 377612 77002 377622
rect 77400 376738 77800 376748
rect 77400 376558 77414 376738
rect 77786 376558 77800 376738
rect 77400 376548 77800 376558
rect 78409 375429 78809 375439
rect 78409 375249 78423 375429
rect 78795 375249 78809 375429
rect 78409 375239 78809 375249
rect 79434 373974 79834 373984
rect 79434 373794 79448 373974
rect 79820 373794 79834 373974
rect 79434 373784 79834 373794
rect 76143 371324 76343 371334
rect 76143 371144 76153 371324
rect 76333 371144 76343 371324
rect 76143 371134 76343 371144
rect 42626 369303 76013 369403
rect 42626 44249 42726 369303
rect 76146 368563 76346 368573
rect 76146 368383 76156 368563
rect 76336 368383 76346 368563
rect 76146 368373 76346 368383
rect 77055 367403 77255 367413
rect 77055 367223 77065 367403
rect 77245 367223 77255 367403
rect 77055 367213 77255 367223
rect 78988 366457 79188 366467
rect 78988 366277 78998 366457
rect 79178 366277 79188 366457
rect 78988 366267 79188 366277
rect 76601 364455 77001 364465
rect 76601 364275 76615 364455
rect 76987 364275 77001 364455
rect 76601 364265 77001 364275
rect 77400 363396 77800 363406
rect 77400 363216 77414 363396
rect 77786 363216 77800 363396
rect 77400 363206 77800 363216
rect 78406 362083 78806 362093
rect 78406 361903 78420 362083
rect 78792 361903 78806 362083
rect 78406 361893 78806 361903
rect 79436 360636 79836 360646
rect 79436 360456 79450 360636
rect 79822 360456 79836 360636
rect 79436 360446 79836 360456
rect 76133 357975 76333 357985
rect 76133 357795 76143 357975
rect 76323 357795 76333 357975
rect 76133 357785 76333 357795
rect 43367 355955 76008 356055
rect 43367 44494 43467 355955
rect 76153 355218 76353 355228
rect 76153 355038 76163 355218
rect 76343 355038 76353 355218
rect 76153 355028 76353 355038
rect 77145 354059 77345 354069
rect 77145 353879 77155 354059
rect 77335 353879 77345 354059
rect 77145 353869 77345 353879
rect 78992 353117 79192 353127
rect 78992 352937 79002 353117
rect 79182 352937 79192 353117
rect 78992 352927 79192 352937
rect 76601 351110 77001 351120
rect 76601 350930 76615 351110
rect 76987 350930 77001 351110
rect 76601 350920 77001 350930
rect 77400 350050 77800 350060
rect 77400 349870 77414 350050
rect 77786 349870 77800 350050
rect 77400 349860 77800 349870
rect 78409 348736 78809 348746
rect 78409 348556 78423 348736
rect 78795 348556 78809 348736
rect 78409 348546 78809 348556
rect 79435 347287 79835 347297
rect 79435 347107 79449 347287
rect 79821 347107 79835 347287
rect 79435 347097 79835 347107
rect 76100 344630 76300 344640
rect 76100 344450 76110 344630
rect 76290 344450 76300 344630
rect 76100 344440 76300 344450
rect 43973 342603 76014 342703
rect 43973 47367 44073 342603
rect 76123 341868 76323 341878
rect 76123 341688 76133 341868
rect 76313 341688 76323 341868
rect 76123 341678 76323 341688
rect 77111 340717 77311 340727
rect 77111 340537 77121 340717
rect 77301 340537 77311 340717
rect 77111 340527 77311 340537
rect 78999 339768 79199 339778
rect 78999 339588 79009 339768
rect 79189 339588 79199 339768
rect 78999 339578 79199 339588
rect 76601 337770 77001 337780
rect 76601 337590 76615 337770
rect 76987 337590 77001 337770
rect 76601 337580 77001 337590
rect 77400 336703 77800 336713
rect 77400 336523 77414 336703
rect 77786 336523 77800 336703
rect 77400 336513 77800 336523
rect 78404 335393 78804 335403
rect 78404 335213 78418 335393
rect 78790 335213 78804 335393
rect 78404 335203 78804 335213
rect 79435 333944 79835 333954
rect 79435 333764 79449 333944
rect 79821 333764 79835 333944
rect 79435 333754 79835 333764
rect 76143 331286 76343 331296
rect 76143 331106 76153 331286
rect 76333 331106 76343 331286
rect 76143 331096 76343 331106
rect 43972 47350 44073 47367
rect 44443 329258 76008 329358
rect 43972 44717 44072 47350
rect 44443 45000 44543 329258
rect 76147 328528 76347 328538
rect 76147 328348 76157 328528
rect 76337 328348 76347 328528
rect 76147 328338 76347 328348
rect 77099 327374 77299 327384
rect 77099 327194 77109 327374
rect 77289 327194 77299 327374
rect 77099 327184 77299 327194
rect 79011 326420 79211 326430
rect 79011 326240 79021 326420
rect 79201 326240 79211 326420
rect 79011 326230 79211 326240
rect 76602 324423 77002 324433
rect 76602 324243 76616 324423
rect 76988 324243 77002 324423
rect 76602 324233 77002 324243
rect 77400 323359 77800 323369
rect 77400 323179 77414 323359
rect 77786 323179 77800 323359
rect 77400 323169 77800 323179
rect 78409 322048 78809 322058
rect 78409 321868 78423 322048
rect 78795 321868 78809 322048
rect 78409 321858 78809 321868
rect 79438 320596 79838 320606
rect 79438 320416 79452 320596
rect 79824 320416 79838 320596
rect 79438 320406 79838 320416
rect 76155 317934 76355 317944
rect 76155 317754 76165 317934
rect 76345 317754 76355 317934
rect 76155 317744 76355 317754
rect 44840 315921 75998 316021
rect 44840 45352 44940 315921
rect 76143 315183 76343 315193
rect 76143 315003 76153 315183
rect 76333 315003 76343 315183
rect 76143 314993 76343 315003
rect 77104 314028 77304 314038
rect 77104 313848 77114 314028
rect 77294 313848 77304 314028
rect 77104 313838 77304 313848
rect 78970 313082 79170 313092
rect 78970 312902 78980 313082
rect 79160 312902 79170 313082
rect 78970 312892 79170 312902
rect 76600 311079 77000 311089
rect 76600 310899 76614 311079
rect 76986 310899 77000 311079
rect 76600 310889 77000 310899
rect 77400 310014 77800 310024
rect 77400 309834 77414 310014
rect 77786 309834 77800 310014
rect 77400 309824 77800 309834
rect 78410 308703 78810 308713
rect 78410 308523 78424 308703
rect 78796 308523 78810 308703
rect 78410 308513 78810 308523
rect 79431 307251 79831 307261
rect 79431 307071 79445 307251
rect 79817 307071 79831 307251
rect 79431 307061 79831 307071
rect 76138 304593 76338 304603
rect 76138 304413 76148 304593
rect 76328 304413 76338 304593
rect 76138 304403 76338 304413
rect 45217 302580 76003 302680
rect 45217 47320 45317 302580
rect 76153 301836 76353 301846
rect 76153 301656 76163 301836
rect 76343 301656 76353 301836
rect 76153 301646 76353 301656
rect 77110 300677 77310 300687
rect 77110 300497 77120 300677
rect 77300 300497 77310 300677
rect 77110 300487 77310 300497
rect 78983 299731 79183 299741
rect 78983 299551 78993 299731
rect 79173 299551 79183 299731
rect 78983 299541 79183 299551
rect 76602 297732 77002 297742
rect 76602 297552 76616 297732
rect 76988 297552 77002 297732
rect 76602 297542 77002 297552
rect 77400 296666 77800 296676
rect 77400 296486 77414 296666
rect 77786 296486 77800 296666
rect 77400 296476 77800 296486
rect 78411 295358 78811 295368
rect 78411 295178 78425 295358
rect 78797 295178 78811 295358
rect 78411 295168 78811 295178
rect 79437 293906 79837 293916
rect 79437 293726 79451 293906
rect 79823 293726 79837 293906
rect 79437 293716 79837 293726
rect 76138 291253 76338 291263
rect 76138 291073 76148 291253
rect 76328 291073 76338 291253
rect 76138 291063 76338 291073
rect 45216 47275 45317 47320
rect 45636 289226 76009 289326
rect 45216 45528 45316 47275
rect 45636 45818 45736 289226
rect 76128 288500 76328 288510
rect 76128 288320 76138 288500
rect 76318 288320 76328 288500
rect 76128 288310 76328 288320
rect 77107 287334 77307 287344
rect 77107 287154 77117 287334
rect 77297 287154 77307 287334
rect 77107 287144 77307 287154
rect 78981 286388 79181 286398
rect 78981 286208 78991 286388
rect 79171 286208 79181 286388
rect 78981 286198 79181 286208
rect 76602 284386 77002 284396
rect 76602 284206 76616 284386
rect 76988 284206 77002 284386
rect 76602 284196 77002 284206
rect 77400 283324 77800 283334
rect 77400 283144 77414 283324
rect 77786 283144 77800 283324
rect 77400 283134 77800 283144
rect 78409 282013 78809 282023
rect 78409 281833 78423 282013
rect 78795 281833 78809 282013
rect 78409 281823 78809 281833
rect 79433 280568 79833 280578
rect 79433 280388 79447 280568
rect 79819 280388 79833 280568
rect 79433 280378 79833 280388
rect 76146 277919 76346 277929
rect 76146 277739 76156 277919
rect 76336 277739 76346 277919
rect 76146 277729 76346 277739
rect 46147 275888 76002 275988
rect 46147 46085 46247 275888
rect 76146 275141 76346 275151
rect 76146 274961 76156 275141
rect 76336 274961 76346 275141
rect 76146 274951 76346 274961
rect 77118 273990 77318 274000
rect 77118 273810 77128 273990
rect 77308 273810 77318 273990
rect 77118 273800 77318 273810
rect 78988 273049 79188 273059
rect 78988 272869 78998 273049
rect 79178 272869 79188 273049
rect 78988 272859 79188 272869
rect 76601 271042 77001 271052
rect 76601 270862 76615 271042
rect 76987 270862 77001 271042
rect 76601 270852 77001 270862
rect 77400 269977 77800 269987
rect 77400 269797 77414 269977
rect 77786 269797 77800 269977
rect 77400 269787 77800 269797
rect 78410 268673 78810 268683
rect 78410 268493 78424 268673
rect 78796 268493 78810 268673
rect 78410 268483 78810 268493
rect 79436 267215 79836 267225
rect 79436 267035 79450 267215
rect 79822 267035 79836 267215
rect 79436 267025 79836 267035
rect 76157 264562 76357 264572
rect 76157 264382 76167 264562
rect 76347 264382 76357 264562
rect 76157 264372 76357 264382
rect 46700 262553 76008 262653
rect 46700 46324 46800 262553
rect 76169 261803 76369 261813
rect 76169 261623 76179 261803
rect 76359 261623 76369 261803
rect 76169 261613 76369 261623
rect 77120 260645 77320 260655
rect 77120 260465 77130 260645
rect 77310 260465 77320 260645
rect 77120 260455 77320 260465
rect 78975 259698 79175 259708
rect 78975 259518 78985 259698
rect 79165 259518 79175 259698
rect 78975 259508 79175 259518
rect 76601 257698 77001 257708
rect 76601 257518 76615 257698
rect 76987 257518 77001 257698
rect 76601 257508 77001 257518
rect 77400 256634 77800 256644
rect 77400 256454 77414 256634
rect 77786 256454 77800 256634
rect 77400 256444 77800 256454
rect 78409 255323 78809 255333
rect 78409 255143 78423 255323
rect 78795 255143 78809 255323
rect 78409 255133 78809 255143
rect 121307 254790 121507 254800
rect 121307 254610 121317 254790
rect 121497 254610 121507 254790
rect 121307 254600 121507 254610
rect 79436 253876 79836 253886
rect 79436 253696 79450 253876
rect 79822 253696 79836 253876
rect 79436 253686 79836 253696
rect 76154 251213 76354 251223
rect 76154 251033 76164 251213
rect 76344 251033 76354 251213
rect 76154 251023 76354 251033
rect 47034 249194 76008 249294
rect 47034 46589 47134 249194
rect 76152 248454 76352 248464
rect 76152 248274 76162 248454
rect 76342 248274 76352 248454
rect 76152 248264 76352 248274
rect 77098 247298 77298 247308
rect 77098 247118 77108 247298
rect 77288 247118 77298 247298
rect 77098 247108 77298 247118
rect 78989 246352 79189 246362
rect 78989 246172 78999 246352
rect 79179 246172 79189 246352
rect 78989 246162 79189 246172
rect 76602 244352 77002 244362
rect 76602 244172 76616 244352
rect 76988 244172 77002 244352
rect 76602 244162 77002 244172
rect 77400 243289 77800 243299
rect 77400 243109 77414 243289
rect 77786 243109 77800 243289
rect 77400 243099 77800 243109
rect 78411 241973 78811 241983
rect 78411 241793 78425 241973
rect 78797 241793 78811 241973
rect 78411 241783 78811 241793
rect 79437 240528 79837 240538
rect 79437 240348 79451 240528
rect 79823 240348 79837 240528
rect 79437 240338 79837 240348
rect 76201 237840 76401 237850
rect 76201 237660 76211 237840
rect 76391 237660 76401 237840
rect 76201 237650 76401 237660
rect 47721 235817 76133 235917
rect 47721 46865 47821 235817
rect 76199 235072 76399 235082
rect 76199 234892 76209 235072
rect 76389 234892 76399 235072
rect 76199 234882 76399 234892
rect 77076 233916 77276 233926
rect 77076 233736 77086 233916
rect 77266 233736 77276 233916
rect 77076 233726 77276 233736
rect 78984 232970 79184 232980
rect 78984 232790 78994 232970
rect 79174 232790 79184 232970
rect 78984 232780 79184 232790
rect 76603 230969 77003 230979
rect 76603 230789 76617 230969
rect 76989 230789 77003 230969
rect 76603 230779 77003 230789
rect 77400 229910 77800 229920
rect 77400 229730 77414 229910
rect 77786 229730 77800 229910
rect 77400 229720 77800 229730
rect 78407 228599 78807 228609
rect 78407 228419 78421 228599
rect 78793 228419 78807 228599
rect 78407 228409 78807 228419
rect 79431 227147 79831 227157
rect 79431 226967 79445 227147
rect 79817 226967 79831 227147
rect 79431 226957 79831 226967
rect 93791 216539 93991 216553
rect 93791 216167 93801 216539
rect 93981 216167 93991 216539
rect 93791 216153 93991 216167
rect 106141 216538 106341 216552
rect 106141 216166 106151 216538
rect 106331 216166 106341 216538
rect 106141 216152 106341 216166
rect 119102 216540 119302 216554
rect 119102 216168 119112 216540
rect 119292 216168 119302 216540
rect 119102 216154 119302 216168
rect 131446 216538 131646 216552
rect 131446 216166 131456 216538
rect 131636 216166 131646 216538
rect 131446 216152 131646 216166
rect 144753 216537 144953 216551
rect 144753 216165 144763 216537
rect 144943 216165 144953 216537
rect 144753 216151 144953 216165
rect 157096 216538 157296 216552
rect 157096 216166 157106 216538
rect 157286 216166 157296 216538
rect 157096 216152 157296 216166
rect 170398 216538 170598 216552
rect 170398 216166 170408 216538
rect 170588 216166 170598 216538
rect 170398 216152 170598 216166
rect 182745 216539 182945 216553
rect 182745 216167 182755 216539
rect 182935 216167 182945 216539
rect 182745 216153 182945 216167
rect 196053 216540 196253 216554
rect 196053 216168 196063 216540
rect 196243 216168 196253 216540
rect 196053 216154 196253 216168
rect 208397 216541 208597 216555
rect 208397 216169 208407 216541
rect 208587 216169 208597 216541
rect 208397 216155 208597 216169
rect 221701 216543 221901 216557
rect 221701 216171 221711 216543
rect 221891 216171 221901 216543
rect 221701 216157 221901 216171
rect 234052 216541 234252 216555
rect 234052 216169 234062 216541
rect 234242 216169 234252 216541
rect 234052 216155 234252 216169
rect 247353 216540 247553 216554
rect 247353 216168 247363 216540
rect 247543 216168 247553 216540
rect 247353 216154 247553 216168
rect 259702 216541 259902 216555
rect 259702 216169 259712 216541
rect 259892 216169 259902 216541
rect 259702 216155 259902 216169
rect 273001 216534 273201 216548
rect 273001 216162 273011 216534
rect 273191 216162 273201 216534
rect 273001 216148 273201 216162
rect 285347 216539 285547 216553
rect 285347 216167 285357 216539
rect 285537 216167 285547 216539
rect 285347 216153 285547 216167
rect 298650 216541 298850 216555
rect 298650 216169 298660 216541
rect 298840 216169 298850 216541
rect 298650 216155 298850 216169
rect 310997 216543 311197 216557
rect 310997 216171 311007 216543
rect 311187 216171 311197 216543
rect 310997 216157 311197 216171
rect 324302 216534 324502 216548
rect 324302 216162 324312 216534
rect 324492 216162 324502 216534
rect 324302 216148 324502 216162
rect 336647 216540 336847 216554
rect 336647 216168 336657 216540
rect 336837 216168 336847 216540
rect 336647 216154 336847 216168
rect 349953 216538 350153 216552
rect 349953 216166 349963 216538
rect 350143 216166 350153 216538
rect 349953 216152 350153 216166
rect 362298 216542 362498 216556
rect 362298 216170 362308 216542
rect 362488 216170 362498 216542
rect 362298 216156 362498 216170
rect 375596 216534 375796 216548
rect 375596 216162 375606 216534
rect 375786 216162 375796 216534
rect 375596 216148 375796 216162
rect 387945 216534 388145 216548
rect 387945 216162 387955 216534
rect 388135 216162 388145 216534
rect 387945 216148 388145 216162
rect 401252 216537 401452 216551
rect 401252 216165 401262 216537
rect 401442 216165 401452 216537
rect 401252 216151 401452 216165
rect 413602 216538 413802 216552
rect 413602 216166 413612 216538
rect 413792 216166 413802 216538
rect 413602 216152 413802 216166
rect 426902 216539 427102 216553
rect 426902 216167 426912 216539
rect 427092 216167 427102 216539
rect 426902 216153 427102 216167
rect 439246 216540 439446 216554
rect 439246 216168 439256 216540
rect 439436 216168 439446 216540
rect 439246 216154 439446 216168
rect 452556 216549 452756 216563
rect 452556 216177 452566 216549
rect 452746 216177 452756 216549
rect 452556 216163 452756 216177
rect 464896 216539 465096 216553
rect 464896 216167 464906 216539
rect 465086 216167 465096 216539
rect 464896 216153 465096 216167
rect 478201 216541 478401 216555
rect 478201 216169 478211 216541
rect 478391 216169 478401 216541
rect 478201 216155 478401 216169
rect 490543 216535 490743 216549
rect 490543 216163 490553 216535
rect 490733 216163 490743 216535
rect 490543 216149 490743 216163
rect 94848 215785 95048 215799
rect 94848 215413 94858 215785
rect 95038 215413 95048 215785
rect 94848 215399 95048 215413
rect 107198 215785 107398 215799
rect 107198 215413 107208 215785
rect 107388 215413 107398 215785
rect 107198 215399 107398 215413
rect 120163 215785 120363 215799
rect 120163 215413 120173 215785
rect 120353 215413 120363 215785
rect 120163 215399 120363 215413
rect 132507 215782 132707 215796
rect 132507 215410 132517 215782
rect 132697 215410 132707 215782
rect 132507 215396 132707 215410
rect 145814 215785 146014 215799
rect 145814 215413 145824 215785
rect 146004 215413 146014 215785
rect 145814 215399 146014 215413
rect 158154 215778 158354 215792
rect 158154 215406 158164 215778
rect 158344 215406 158354 215778
rect 158154 215392 158354 215406
rect 171464 215784 171664 215798
rect 171464 215412 171474 215784
rect 171654 215412 171664 215784
rect 171464 215398 171664 215412
rect 183807 215785 184007 215799
rect 183807 215413 183817 215785
rect 183997 215413 184007 215785
rect 183807 215399 184007 215413
rect 197110 215786 197310 215800
rect 197110 215414 197120 215786
rect 197300 215414 197310 215786
rect 197110 215400 197310 215414
rect 209458 215786 209658 215800
rect 209458 215414 209468 215786
rect 209648 215414 209658 215786
rect 209458 215400 209658 215414
rect 222764 215786 222964 215800
rect 222764 215414 222774 215786
rect 222954 215414 222964 215786
rect 222764 215400 222964 215414
rect 235107 215786 235307 215800
rect 235107 215414 235117 215786
rect 235297 215414 235307 215786
rect 235107 215400 235307 215414
rect 248409 215785 248609 215799
rect 248409 215413 248419 215785
rect 248599 215413 248609 215785
rect 248409 215399 248609 215413
rect 260760 215786 260960 215800
rect 260760 215414 260770 215786
rect 260950 215414 260960 215786
rect 260760 215400 260960 215414
rect 274061 215784 274261 215798
rect 274061 215412 274071 215784
rect 274251 215412 274261 215784
rect 274061 215398 274261 215412
rect 286405 215784 286605 215798
rect 286405 215412 286415 215784
rect 286595 215412 286605 215784
rect 286405 215398 286605 215412
rect 299709 215786 299909 215800
rect 299709 215414 299719 215786
rect 299899 215414 299909 215786
rect 299709 215400 299909 215414
rect 312056 215786 312256 215800
rect 312056 215414 312066 215786
rect 312246 215414 312256 215786
rect 312056 215400 312256 215414
rect 325361 215784 325561 215798
rect 325361 215412 325371 215784
rect 325551 215412 325561 215784
rect 325361 215398 325561 215412
rect 337706 215781 337906 215795
rect 337706 215409 337716 215781
rect 337896 215409 337906 215781
rect 337706 215395 337906 215409
rect 351008 215784 351208 215798
rect 351008 215412 351018 215784
rect 351198 215412 351208 215784
rect 351008 215398 351208 215412
rect 363357 215784 363557 215798
rect 363357 215412 363367 215784
rect 363547 215412 363557 215784
rect 363357 215398 363557 215412
rect 376662 215781 376862 215795
rect 376662 215409 376672 215781
rect 376852 215409 376862 215781
rect 376662 215395 376862 215409
rect 389004 215787 389204 215801
rect 389004 215415 389014 215787
rect 389194 215415 389204 215787
rect 389004 215401 389204 215415
rect 402311 215783 402511 215797
rect 402311 215411 402321 215783
rect 402501 215411 402511 215783
rect 402311 215397 402511 215411
rect 414658 215781 414858 215795
rect 414658 215409 414668 215781
rect 414848 215409 414858 215781
rect 414658 215395 414858 215409
rect 427961 215788 428161 215802
rect 427961 215416 427971 215788
rect 428151 215416 428161 215788
rect 427961 215402 428161 215416
rect 440306 215782 440506 215796
rect 440306 215410 440316 215782
rect 440496 215410 440506 215782
rect 440306 215396 440506 215410
rect 453612 215788 453812 215802
rect 453612 215416 453622 215788
rect 453802 215416 453812 215788
rect 453612 215402 453812 215416
rect 465958 215786 466158 215800
rect 465958 215414 465968 215786
rect 466148 215414 466158 215786
rect 465958 215400 466158 215414
rect 479259 215784 479459 215798
rect 479259 215412 479269 215784
rect 479449 215412 479459 215784
rect 479259 215398 479459 215412
rect 491606 215784 491806 215798
rect 491606 215412 491616 215784
rect 491796 215412 491806 215784
rect 491606 215398 491806 215412
rect 257695 215290 257895 215300
rect 232046 215275 232246 215285
rect 117109 215263 117309 215273
rect 91790 215250 91990 215260
rect 91790 215070 91800 215250
rect 91980 215070 91990 215250
rect 91790 215060 91990 215070
rect 104135 215241 104335 215251
rect 104135 215061 104145 215241
rect 104325 215061 104335 215241
rect 117109 215083 117119 215263
rect 117299 215083 117309 215263
rect 194044 215263 194244 215273
rect 155099 215247 155299 215257
rect 142759 215217 142959 215227
rect 117109 215073 117309 215083
rect 129444 215201 129644 215211
rect 104135 215051 104335 215061
rect 129444 215021 129454 215201
rect 129634 215021 129644 215201
rect 142759 215037 142769 215217
rect 142949 215037 142959 215217
rect 155099 215067 155109 215247
rect 155289 215067 155299 215247
rect 180755 215235 180955 215245
rect 155099 215057 155299 215067
rect 168401 215204 168601 215214
rect 142759 215027 142959 215037
rect 129444 215011 129644 215021
rect 168401 215024 168411 215204
rect 168591 215024 168601 215204
rect 180755 215055 180765 215235
rect 180945 215055 180955 215235
rect 194044 215083 194054 215263
rect 194234 215083 194244 215263
rect 194044 215073 194244 215083
rect 206402 215241 206602 215251
rect 180755 215045 180955 215055
rect 206402 215061 206412 215241
rect 206592 215061 206602 215241
rect 206402 215051 206602 215061
rect 219699 215240 219899 215250
rect 219699 215060 219709 215240
rect 219889 215060 219899 215240
rect 232046 215095 232056 215275
rect 232236 215095 232246 215275
rect 232046 215085 232246 215095
rect 245350 215259 245550 215269
rect 245350 215079 245360 215259
rect 245540 215079 245550 215259
rect 257695 215110 257705 215290
rect 257885 215110 257895 215290
rect 257695 215100 257895 215110
rect 271004 215271 271204 215281
rect 271004 215091 271014 215271
rect 271194 215091 271204 215271
rect 271004 215081 271204 215091
rect 283347 215253 283547 215263
rect 245350 215069 245550 215079
rect 283347 215073 283357 215253
rect 283537 215073 283547 215253
rect 283347 215063 283547 215073
rect 296650 215249 296850 215259
rect 296650 215069 296660 215249
rect 296840 215069 296850 215249
rect 219699 215050 219899 215060
rect 296650 215059 296850 215069
rect 308994 215256 309194 215266
rect 308994 215076 309004 215256
rect 309184 215076 309194 215256
rect 334645 215263 334845 215273
rect 308994 215066 309194 215076
rect 322301 215233 322501 215243
rect 322301 215053 322311 215233
rect 322491 215053 322501 215233
rect 334645 215083 334655 215263
rect 334835 215083 334845 215263
rect 385945 215264 386145 215274
rect 360295 215245 360495 215255
rect 334645 215073 334845 215083
rect 347951 215233 348151 215243
rect 322301 215043 322501 215053
rect 347951 215053 347961 215233
rect 348141 215053 348151 215233
rect 360295 215065 360305 215245
rect 360485 215065 360495 215245
rect 360295 215055 360495 215065
rect 373600 215237 373800 215247
rect 373600 215057 373610 215237
rect 373790 215057 373800 215237
rect 385945 215084 385955 215264
rect 386135 215084 386145 215264
rect 385945 215074 386145 215084
rect 399250 215263 399450 215273
rect 399250 215083 399260 215263
rect 399440 215083 399450 215263
rect 437247 215250 437447 215260
rect 399250 215073 399450 215083
rect 411599 215229 411799 215239
rect 347951 215043 348151 215053
rect 373600 215047 373800 215057
rect 411599 215049 411609 215229
rect 411789 215049 411799 215229
rect 411599 215039 411799 215049
rect 424899 215232 425099 215242
rect 424899 215052 424909 215232
rect 425089 215052 425099 215232
rect 437247 215070 437257 215250
rect 437437 215070 437447 215250
rect 437247 215060 437447 215070
rect 450543 215250 450743 215260
rect 450543 215070 450553 215250
rect 450733 215070 450743 215250
rect 450543 215060 450743 215070
rect 462894 215237 463094 215247
rect 424899 215042 425099 215052
rect 462894 215057 462904 215237
rect 463084 215057 463094 215237
rect 488547 215243 488747 215253
rect 462894 215047 463094 215057
rect 476206 215225 476406 215235
rect 476206 215045 476216 215225
rect 476396 215045 476406 215225
rect 488547 215063 488557 215243
rect 488737 215063 488747 215243
rect 488547 215053 488747 215063
rect 476206 215035 476406 215045
rect 168401 215014 168601 215024
rect 96165 214904 96365 214918
rect 96165 214532 96175 214904
rect 96355 214532 96365 214904
rect 96165 214518 96365 214532
rect 108508 214907 108708 214921
rect 108508 214535 108518 214907
rect 108698 214535 108708 214907
rect 108508 214521 108708 214535
rect 121474 214901 121674 214915
rect 121474 214529 121484 214901
rect 121664 214529 121674 214901
rect 121474 214515 121674 214529
rect 133818 214903 134018 214917
rect 133818 214531 133828 214903
rect 134008 214531 134018 214903
rect 133818 214517 134018 214531
rect 147122 214903 147322 214917
rect 147122 214531 147132 214903
rect 147312 214531 147322 214903
rect 147122 214517 147322 214531
rect 159470 214906 159670 214920
rect 159470 214534 159480 214906
rect 159660 214534 159670 214906
rect 159470 214520 159670 214534
rect 172774 214904 172974 214918
rect 172774 214532 172784 214904
rect 172964 214532 172974 214904
rect 172774 214518 172974 214532
rect 185121 214904 185321 214918
rect 185121 214532 185131 214904
rect 185311 214532 185321 214904
rect 185121 214518 185321 214532
rect 198422 214902 198622 214916
rect 198422 214530 198432 214902
rect 198612 214530 198622 214902
rect 198422 214516 198622 214530
rect 210771 214903 210971 214917
rect 210771 214531 210781 214903
rect 210961 214531 210971 214903
rect 210771 214517 210971 214531
rect 224078 214906 224278 214920
rect 224078 214534 224088 214906
rect 224268 214534 224278 214906
rect 224078 214520 224278 214534
rect 236418 214904 236618 214918
rect 236418 214532 236428 214904
rect 236608 214532 236618 214904
rect 236418 214518 236618 214532
rect 249722 214901 249922 214915
rect 249722 214529 249732 214901
rect 249912 214529 249922 214901
rect 249722 214515 249922 214529
rect 262070 214905 262270 214919
rect 262070 214533 262080 214905
rect 262260 214533 262270 214905
rect 262070 214519 262270 214533
rect 275373 214903 275573 214917
rect 275373 214531 275383 214903
rect 275563 214531 275573 214903
rect 275373 214517 275573 214531
rect 287721 214903 287921 214917
rect 287721 214531 287731 214903
rect 287911 214531 287921 214903
rect 287721 214517 287921 214531
rect 301030 214906 301230 214920
rect 301030 214534 301040 214906
rect 301220 214534 301230 214906
rect 301030 214520 301230 214534
rect 313368 214904 313568 214918
rect 313368 214532 313378 214904
rect 313558 214532 313568 214904
rect 313368 214518 313568 214532
rect 326673 214903 326873 214917
rect 326673 214531 326683 214903
rect 326863 214531 326873 214903
rect 326673 214517 326873 214531
rect 339018 214904 339218 214918
rect 339018 214532 339028 214904
rect 339208 214532 339218 214904
rect 339018 214518 339218 214532
rect 352324 214901 352524 214915
rect 352324 214529 352334 214901
rect 352514 214529 352524 214901
rect 352324 214515 352524 214529
rect 364669 214904 364869 214918
rect 364669 214532 364679 214904
rect 364859 214532 364869 214904
rect 364669 214518 364869 214532
rect 377974 214904 378174 214918
rect 377974 214532 377984 214904
rect 378164 214532 378174 214904
rect 377974 214518 378174 214532
rect 390321 214902 390521 214916
rect 390321 214530 390331 214902
rect 390511 214530 390521 214902
rect 390321 214516 390521 214530
rect 403614 214894 403814 214908
rect 403614 214522 403624 214894
rect 403804 214522 403814 214894
rect 403614 214508 403814 214522
rect 415966 214898 416166 214912
rect 415966 214526 415976 214898
rect 416156 214526 416166 214898
rect 415966 214512 416166 214526
rect 429276 214901 429476 214915
rect 429276 214529 429286 214901
rect 429466 214529 429476 214901
rect 429276 214515 429476 214529
rect 441618 214904 441818 214918
rect 441618 214532 441628 214904
rect 441808 214532 441818 214904
rect 441618 214518 441818 214532
rect 454924 214907 455124 214921
rect 454924 214535 454934 214907
rect 455114 214535 455124 214907
rect 454924 214521 455124 214535
rect 467268 214902 467468 214916
rect 467268 214530 467278 214902
rect 467458 214530 467468 214902
rect 467268 214516 467468 214530
rect 480569 214901 480769 214915
rect 480569 214529 480579 214901
rect 480759 214529 480769 214901
rect 480569 214515 480769 214529
rect 492922 214902 493122 214916
rect 492922 214530 492932 214902
rect 493112 214530 493122 214902
rect 492922 214516 493122 214530
rect 97613 214115 97813 214129
rect 97613 213743 97623 214115
rect 97803 213743 97813 214115
rect 97613 213729 97813 213743
rect 109971 214111 110171 214125
rect 109971 213739 109981 214111
rect 110161 213739 110171 214111
rect 109971 213725 110171 213739
rect 122925 214116 123125 214130
rect 122925 213744 122935 214116
rect 123115 213744 123125 214116
rect 122925 213730 123125 213744
rect 135288 214113 135488 214127
rect 135288 213741 135298 214113
rect 135478 213741 135488 214113
rect 135288 213727 135488 213741
rect 148581 214105 148781 214119
rect 148581 213733 148591 214105
rect 148771 213733 148781 214105
rect 148581 213719 148781 213733
rect 160921 214105 161121 214119
rect 160921 213733 160931 214105
rect 161111 213733 161121 214105
rect 160921 213719 161121 213733
rect 174225 214111 174425 214125
rect 174225 213739 174235 214111
rect 174415 213739 174425 214111
rect 174225 213725 174425 213739
rect 186585 214123 186785 214137
rect 186585 213751 186595 214123
rect 186775 213751 186785 214123
rect 212226 214119 212426 214133
rect 186585 213737 186785 213751
rect 199877 214105 200077 214119
rect 199877 213733 199887 214105
rect 200067 213733 200077 214105
rect 212226 213747 212236 214119
rect 212416 213747 212426 214119
rect 212226 213733 212426 213747
rect 225532 214113 225732 214127
rect 225532 213741 225542 214113
rect 225722 213741 225732 214113
rect 199877 213719 200077 213733
rect 225532 213727 225732 213741
rect 237886 214115 238086 214129
rect 237886 213743 237896 214115
rect 238076 213743 238086 214115
rect 237886 213729 238086 213743
rect 251189 214116 251389 214130
rect 251189 213744 251199 214116
rect 251379 213744 251389 214116
rect 251189 213730 251389 213744
rect 263531 214120 263731 214134
rect 263531 213748 263541 214120
rect 263721 213748 263731 214120
rect 263531 213734 263731 213748
rect 276838 214111 277038 214125
rect 276838 213739 276848 214111
rect 277028 213739 277038 214111
rect 276838 213725 277038 213739
rect 289167 214110 289367 214124
rect 289167 213738 289177 214110
rect 289357 213738 289367 214110
rect 289167 213724 289367 213738
rect 302486 214113 302686 214127
rect 302486 213741 302496 214113
rect 302676 213741 302686 214113
rect 302486 213727 302686 213741
rect 314825 214116 315025 214130
rect 314825 213744 314835 214116
rect 315015 213744 315025 214116
rect 314825 213730 315025 213744
rect 328123 214116 328323 214130
rect 328123 213744 328133 214116
rect 328313 213744 328323 214116
rect 328123 213730 328323 213744
rect 340473 214117 340673 214131
rect 340473 213745 340483 214117
rect 340663 213745 340673 214117
rect 340473 213731 340673 213745
rect 353782 214113 353982 214127
rect 353782 213741 353792 214113
rect 353972 213741 353982 214113
rect 353782 213727 353982 213741
rect 366116 214118 366316 214132
rect 366116 213746 366126 214118
rect 366306 213746 366316 214118
rect 366116 213732 366316 213746
rect 379434 214117 379634 214131
rect 379434 213745 379444 214117
rect 379624 213745 379634 214117
rect 379434 213731 379634 213745
rect 391768 214114 391968 214128
rect 391768 213742 391778 214114
rect 391958 213742 391968 214114
rect 391768 213728 391968 213742
rect 405079 214110 405279 214124
rect 405079 213738 405089 214110
rect 405269 213738 405279 214110
rect 405079 213724 405279 213738
rect 417427 214120 417627 214134
rect 417427 213748 417437 214120
rect 417617 213748 417627 214120
rect 417427 213734 417627 213748
rect 430742 214119 430942 214133
rect 430742 213747 430752 214119
rect 430932 213747 430942 214119
rect 430742 213733 430942 213747
rect 443078 214113 443278 214127
rect 443078 213741 443088 214113
rect 443268 213741 443278 214113
rect 443078 213727 443278 213741
rect 456383 214113 456583 214127
rect 456383 213741 456393 214113
rect 456573 213741 456583 214113
rect 456383 213727 456583 213741
rect 468736 214119 468936 214133
rect 468736 213747 468746 214119
rect 468926 213747 468936 214119
rect 468736 213733 468936 213747
rect 482038 214113 482238 214127
rect 482038 213741 482048 214113
rect 482228 213741 482238 214113
rect 482038 213727 482238 213741
rect 494373 214114 494573 214128
rect 494373 213742 494383 214114
rect 494563 213742 494573 214114
rect 494373 213728 494573 213742
rect 436200 213529 436600 213543
rect 90843 213445 91043 213455
rect 90843 213265 90853 213445
rect 91033 213265 91043 213445
rect 90843 213255 91043 213265
rect 103193 213443 103393 213453
rect 103193 213263 103203 213443
rect 103383 213263 103393 213443
rect 103193 213253 103393 213263
rect 116153 213444 116353 213454
rect 116153 213264 116163 213444
rect 116343 213264 116353 213444
rect 347002 213441 347202 213451
rect 154145 213428 154345 213438
rect 116153 213254 116353 213264
rect 128496 213403 128696 213413
rect 128496 213223 128506 213403
rect 128686 213223 128696 213403
rect 128496 213213 128696 213223
rect 141801 213363 142001 213373
rect 141801 213183 141811 213363
rect 141991 213183 142001 213363
rect 154145 213248 154155 213428
rect 154335 213248 154345 213428
rect 179800 213423 180000 213433
rect 205446 213429 205646 213439
rect 154145 213238 154345 213248
rect 167456 213389 167656 213399
rect 167456 213209 167466 213389
rect 167646 213209 167656 213389
rect 179800 213243 179810 213423
rect 179990 213243 180000 213423
rect 179800 213233 180000 213243
rect 193110 213415 193310 213425
rect 193110 213235 193120 213415
rect 193300 213235 193310 213415
rect 205446 213249 205456 213429
rect 205636 213249 205646 213429
rect 205446 213239 205646 213249
rect 218751 213430 218951 213440
rect 218751 213250 218761 213430
rect 218941 213250 218951 213430
rect 256749 213427 256949 213437
rect 218751 213240 218951 213250
rect 231101 213417 231301 213427
rect 193110 213225 193310 213235
rect 231101 213237 231111 213417
rect 231291 213237 231301 213417
rect 231101 213227 231301 213237
rect 244400 213407 244600 213417
rect 244400 213227 244410 213407
rect 244590 213227 244600 213407
rect 256749 213247 256759 213427
rect 256939 213247 256949 213427
rect 256749 213237 256949 213247
rect 270058 213408 270258 213418
rect 321351 213417 321551 213427
rect 244400 213217 244600 213227
rect 270058 213228 270068 213408
rect 270248 213228 270258 213408
rect 295705 213400 295905 213410
rect 270058 213218 270258 213228
rect 282402 213385 282602 213395
rect 167456 213199 167656 213209
rect 282402 213205 282412 213385
rect 282592 213205 282602 213385
rect 295705 213220 295715 213400
rect 295895 213220 295905 213400
rect 295705 213210 295905 213220
rect 308053 213358 308253 213368
rect 282402 213195 282602 213205
rect 141801 213173 142001 213183
rect 308053 213178 308063 213358
rect 308243 213178 308253 213358
rect 321351 213237 321361 213417
rect 321541 213237 321551 213417
rect 321351 213227 321551 213237
rect 333696 213374 333896 213384
rect 333696 213194 333706 213374
rect 333886 213194 333896 213374
rect 347002 213261 347012 213441
rect 347192 213261 347202 213441
rect 372654 213441 372854 213451
rect 347002 213251 347202 213261
rect 359351 213429 359551 213439
rect 359351 213249 359361 213429
rect 359541 213249 359551 213429
rect 372654 213261 372664 213441
rect 372844 213261 372854 213441
rect 372654 213251 372854 213261
rect 385001 213442 385201 213452
rect 385001 213262 385011 213442
rect 385191 213262 385201 213442
rect 385001 213252 385201 213262
rect 398298 213437 398498 213447
rect 398298 213257 398308 213437
rect 398488 213257 398498 213437
rect 359351 213239 359551 213249
rect 398298 213247 398498 213257
rect 410646 213437 410846 213447
rect 410646 213257 410656 213437
rect 410836 213257 410846 213437
rect 410646 213247 410846 213257
rect 423955 213440 424155 213450
rect 423955 213260 423965 213440
rect 424145 213260 424155 213440
rect 423955 213250 424155 213260
rect 333696 213184 333896 213194
rect 308053 213168 308253 213178
rect 436200 213157 436214 213529
rect 436586 213157 436600 213529
rect 449605 213433 449805 213443
rect 449605 213253 449615 213433
rect 449795 213253 449805 213433
rect 449605 213243 449805 213253
rect 461953 213431 462153 213441
rect 461953 213251 461963 213431
rect 462143 213251 462153 213431
rect 461953 213241 462153 213251
rect 475250 213426 475450 213436
rect 475250 213246 475260 213426
rect 475440 213246 475450 213426
rect 475250 213236 475450 213246
rect 487598 213400 487798 213410
rect 487598 213220 487608 213400
rect 487788 213220 487798 213400
rect 487598 213210 487798 213220
rect 436200 213143 436600 213157
rect 86929 212784 87129 212794
rect 86929 212604 86939 212784
rect 87119 212604 87129 212784
rect 115001 212793 115201 212803
rect 112234 212768 112434 212778
rect 86929 212594 87129 212604
rect 89691 212753 89891 212763
rect 89691 212573 89701 212753
rect 89881 212573 89891 212753
rect 102047 212758 102247 212768
rect 89691 212563 89891 212573
rect 99274 212733 99474 212743
rect 99274 212553 99284 212733
rect 99464 212553 99474 212733
rect 102047 212578 102057 212758
rect 102237 212578 102247 212758
rect 112234 212588 112244 212768
rect 112424 212588 112434 212768
rect 115001 212613 115011 212793
rect 115191 212613 115201 212793
rect 332544 212788 332744 212798
rect 115001 212603 115201 212613
rect 124573 212758 124773 212768
rect 140651 212765 140851 212775
rect 112234 212578 112434 212588
rect 124573 212578 124583 212758
rect 124763 212578 124773 212758
rect 102047 212568 102247 212578
rect 124573 212568 124773 212578
rect 127346 212749 127546 212759
rect 127346 212569 127356 212749
rect 127536 212569 127546 212749
rect 127346 212559 127546 212569
rect 137889 212745 138089 212755
rect 137889 212565 137899 212745
rect 138079 212565 138089 212745
rect 140651 212585 140661 212765
rect 140841 212585 140851 212765
rect 214834 212767 215034 212777
rect 201526 212747 201726 212757
rect 152989 212722 153189 212732
rect 140651 212575 140851 212585
rect 150231 212706 150431 212716
rect 137889 212555 138089 212565
rect 99274 212543 99474 212553
rect 150231 212526 150241 212706
rect 150421 212526 150431 212706
rect 152989 212542 152999 212722
rect 153179 212542 153189 212722
rect 152989 212532 153189 212542
rect 163531 212723 163731 212733
rect 163531 212543 163541 212723
rect 163721 212543 163731 212723
rect 175881 212730 176081 212740
rect 163531 212533 163731 212543
rect 166302 212711 166502 212721
rect 150231 212516 150431 212526
rect 166302 212531 166312 212711
rect 166492 212531 166502 212711
rect 175881 212550 175891 212730
rect 176071 212550 176081 212730
rect 189185 212737 189385 212747
rect 175881 212540 176081 212550
rect 178642 212711 178842 212721
rect 166302 212521 166502 212531
rect 178642 212531 178652 212711
rect 178832 212531 178842 212711
rect 189185 212557 189195 212737
rect 189375 212557 189385 212737
rect 189185 212547 189385 212557
rect 191952 212737 192152 212747
rect 191952 212557 191962 212737
rect 192142 212557 192152 212737
rect 201526 212567 201536 212747
rect 201716 212567 201726 212747
rect 201526 212557 201726 212567
rect 204292 212725 204492 212735
rect 191952 212547 192152 212557
rect 204292 212545 204302 212725
rect 204482 212545 204492 212725
rect 214834 212587 214844 212767
rect 215024 212587 215034 212767
rect 214834 212577 215034 212587
rect 217598 212763 217798 212773
rect 217598 212583 217608 212763
rect 217788 212583 217798 212763
rect 217598 212573 217798 212583
rect 227185 212756 227385 212766
rect 227185 212576 227195 212756
rect 227375 212576 227385 212756
rect 240486 212755 240686 212765
rect 227185 212566 227385 212576
rect 229944 212734 230144 212744
rect 204292 212535 204492 212545
rect 229944 212554 229954 212734
rect 230134 212554 230144 212734
rect 240486 212575 240496 212755
rect 240676 212575 240686 212755
rect 240486 212565 240686 212575
rect 243247 212764 243447 212774
rect 243247 212584 243257 212764
rect 243437 212584 243447 212764
rect 243247 212574 243447 212584
rect 252832 212745 253032 212755
rect 252832 212565 252842 212745
rect 253022 212565 253032 212745
rect 252832 212555 253032 212565
rect 255592 212745 255792 212755
rect 329781 212753 329981 212763
rect 255592 212565 255602 212745
rect 255782 212565 255792 212745
rect 281245 212736 281445 212746
rect 278477 212726 278677 212736
rect 268900 212695 269100 212705
rect 255592 212555 255792 212565
rect 266133 212661 266333 212671
rect 229944 212544 230144 212554
rect 178642 212521 178842 212531
rect 266133 212481 266143 212661
rect 266323 212481 266333 212661
rect 268900 212515 268910 212695
rect 269090 212515 269100 212695
rect 278477 212546 278487 212726
rect 278667 212546 278677 212726
rect 281245 212556 281255 212736
rect 281435 212556 281445 212736
rect 317440 212726 317640 212736
rect 304137 212711 304337 212721
rect 294548 212691 294748 212701
rect 281245 212546 281445 212556
rect 291785 212670 291985 212680
rect 278477 212536 278677 212546
rect 268900 212505 269100 212515
rect 266133 212471 266333 212481
rect 291785 212490 291795 212670
rect 291975 212490 291985 212670
rect 294548 212511 294558 212691
rect 294738 212511 294748 212691
rect 304137 212531 304147 212711
rect 304327 212531 304337 212711
rect 304137 212521 304337 212531
rect 306901 212706 307101 212716
rect 306901 212526 306911 212706
rect 307091 212526 307101 212706
rect 317440 212546 317450 212726
rect 317630 212546 317640 212726
rect 317440 212536 317640 212546
rect 320198 212726 320398 212736
rect 320198 212546 320208 212726
rect 320388 212546 320398 212726
rect 329781 212573 329791 212753
rect 329971 212573 329981 212753
rect 332544 212608 332554 212788
rect 332734 212608 332744 212788
rect 383846 212772 384046 212782
rect 381081 212753 381281 212763
rect 358194 212739 358394 212749
rect 332544 212598 332744 212608
rect 343087 212724 343287 212734
rect 329781 212563 329981 212573
rect 320198 212536 320398 212546
rect 343087 212544 343097 212724
rect 343277 212544 343287 212724
rect 343087 212534 343287 212544
rect 345849 212729 346049 212739
rect 345849 212549 345859 212729
rect 346039 212549 346049 212729
rect 345849 212539 346049 212549
rect 355428 212720 355628 212730
rect 355428 212540 355438 212720
rect 355618 212540 355628 212720
rect 358194 212559 358204 212739
rect 358384 212559 358394 212739
rect 371499 212730 371699 212740
rect 358194 212549 358394 212559
rect 368737 212706 368937 212716
rect 355428 212530 355628 212540
rect 306901 212516 307101 212526
rect 368737 212526 368747 212706
rect 368927 212526 368937 212706
rect 371499 212550 371509 212730
rect 371689 212550 371699 212730
rect 381081 212573 381091 212753
rect 381271 212573 381281 212753
rect 383846 212592 383856 212772
rect 384036 212592 384046 212772
rect 397149 212767 397349 212777
rect 422800 212776 423000 212786
rect 383846 212582 384046 212592
rect 394388 212717 394588 212727
rect 381081 212563 381281 212573
rect 371499 212540 371699 212550
rect 394388 212537 394398 212717
rect 394578 212537 394588 212717
rect 397149 212587 397159 212767
rect 397339 212587 397349 212767
rect 409496 212753 409696 212763
rect 397149 212577 397349 212587
rect 406727 212733 406927 212743
rect 406727 212553 406737 212733
rect 406917 212553 406927 212733
rect 409496 212573 409506 212753
rect 409686 212573 409696 212753
rect 409496 212563 409696 212573
rect 420037 212758 420237 212768
rect 420037 212578 420047 212758
rect 420227 212578 420237 212758
rect 422800 212596 422810 212776
rect 422990 212596 423000 212776
rect 422800 212586 423000 212596
rect 432386 212773 432586 212783
rect 432386 212593 432396 212773
rect 432576 212593 432586 212773
rect 432386 212583 432586 212593
rect 435145 212745 435345 212755
rect 420037 212568 420237 212578
rect 435145 212565 435155 212745
rect 435335 212565 435345 212745
rect 448449 212744 448649 212754
rect 435145 212555 435345 212565
rect 445681 212690 445881 212700
rect 406727 212543 406927 212553
rect 394388 212527 394588 212537
rect 368737 212516 368937 212526
rect 294548 212501 294748 212511
rect 445681 212510 445691 212690
rect 445871 212510 445881 212690
rect 448449 212564 448459 212744
rect 448639 212564 448649 212744
rect 460793 212737 460993 212747
rect 448449 212554 448649 212564
rect 458031 212705 458231 212715
rect 458031 212525 458041 212705
rect 458221 212525 458231 212705
rect 460793 212557 460803 212737
rect 460983 212557 460993 212737
rect 486447 212741 486647 212751
rect 474100 212713 474300 212723
rect 460793 212547 460993 212557
rect 471328 212659 471528 212669
rect 458031 212515 458231 212525
rect 445681 212500 445881 212510
rect 291785 212480 291985 212490
rect 471328 212479 471338 212659
rect 471518 212479 471528 212659
rect 474100 212533 474110 212713
rect 474290 212533 474300 212713
rect 474100 212523 474300 212533
rect 483684 212671 483884 212681
rect 483684 212491 483694 212671
rect 483874 212491 483884 212671
rect 486447 212561 486457 212741
rect 486637 212561 486647 212741
rect 486447 212551 486647 212561
rect 483684 212481 483884 212491
rect 471328 212469 471528 212479
rect 87881 211604 87981 212279
rect 57717 211504 87981 211604
rect 57717 61817 57817 211504
rect 113186 210948 113286 212295
rect 57990 210848 113286 210948
rect 57990 62551 58090 210848
rect 138854 210142 138954 212327
rect 58330 210042 138954 210142
rect 58330 63378 58430 210042
rect 164497 209449 164597 212304
rect 59385 209349 164597 209449
rect 59385 64222 59485 209349
rect 190149 208571 190249 212343
rect 60453 208471 190249 208571
rect 60453 65376 60553 208471
rect 215797 207826 215897 212336
rect 61307 207726 215897 207826
rect 61307 66672 61407 207726
rect 241446 207154 241546 212344
rect 61869 207054 241546 207154
rect 61869 67306 61969 207054
rect 267100 204457 267200 212333
rect 63249 204357 267200 204457
rect 63249 69658 63349 204357
rect 292738 203747 292838 212332
rect 64105 203647 292838 203747
rect 64105 70545 64205 203647
rect 318401 201530 318501 212337
rect 66302 201430 318501 201530
rect 66302 71921 66402 201430
rect 344038 200319 344138 212335
rect 67891 200219 344138 200319
rect 67891 73266 67991 200219
rect 369693 199242 369793 212342
rect 68994 199142 369793 199242
rect 68994 74343 69094 199142
rect 395339 197097 395439 212339
rect 70189 196997 395439 197097
rect 70189 75161 70289 196997
rect 420990 196045 421090 212338
rect 73133 195945 421090 196045
rect 73133 76808 73233 195945
rect 446638 195150 446738 212337
rect 74184 195050 446738 195150
rect 74184 77859 74284 195050
rect 472290 193724 472390 212338
rect 75185 193624 472390 193724
rect 75185 78919 75285 193624
rect 75185 78895 292684 78919
rect 75185 78843 292516 78895
rect 292568 78843 292684 78895
rect 75185 78819 292684 78843
rect 74184 77835 289130 77859
rect 74184 77783 288955 77835
rect 289007 77783 289130 77835
rect 74184 77759 289130 77783
rect 73133 76784 285571 76808
rect 73133 76732 285422 76784
rect 285474 76732 285571 76784
rect 73133 76708 285571 76732
rect 70189 75137 282030 75161
rect 70189 75085 281872 75137
rect 281924 75085 282030 75137
rect 70189 75061 282030 75085
rect 68994 74319 278491 74343
rect 68994 74267 278312 74319
rect 278364 74267 278491 74319
rect 68994 74243 278491 74267
rect 67891 73242 274969 73266
rect 67891 73190 274773 73242
rect 274825 73190 274969 73242
rect 67891 73166 274969 73190
rect 66302 71897 271447 71921
rect 66302 71845 271233 71897
rect 271285 71845 271447 71897
rect 66302 71821 271447 71845
rect 64105 70521 267849 70545
rect 64105 70469 267693 70521
rect 267745 70469 267849 70521
rect 64105 70445 267849 70469
rect 63249 69634 264326 69658
rect 63249 69582 264145 69634
rect 264197 69582 264326 69634
rect 63249 69558 264326 69582
rect 61869 67282 260747 67306
rect 61869 67230 260593 67282
rect 260645 67230 260747 67282
rect 61869 67206 260747 67230
rect 61307 66648 257229 66672
rect 61307 66596 257049 66648
rect 257101 66596 257229 66648
rect 61307 66572 257229 66596
rect 60453 65352 253682 65376
rect 60453 65300 253511 65352
rect 253563 65300 253682 65352
rect 60453 65276 253682 65300
rect 59385 64198 250131 64222
rect 59385 64146 249945 64198
rect 249997 64146 250131 64198
rect 59385 64122 250131 64146
rect 246360 63378 246460 63379
rect 58330 63355 246605 63378
rect 58330 63303 246384 63355
rect 246436 63303 246605 63355
rect 58330 63278 246605 63303
rect 57990 62527 243038 62551
rect 57990 62475 242866 62527
rect 242918 62475 243038 62527
rect 57990 62451 243038 62475
rect 57717 61793 239537 61817
rect 57717 61741 239313 61793
rect 239365 61741 239537 61793
rect 57717 61717 239537 61741
rect 47721 46841 179167 46865
rect 47721 46789 179041 46841
rect 179093 46789 179167 46841
rect 47721 46765 179167 46789
rect 47034 46565 175620 46589
rect 47034 46513 175484 46565
rect 175536 46513 175620 46565
rect 47034 46489 175620 46513
rect 46700 46300 172089 46324
rect 46700 46248 171955 46300
rect 172007 46248 172089 46300
rect 46700 46224 172089 46248
rect 46147 46061 168542 46085
rect 46147 46009 168401 46061
rect 168453 46009 168542 46061
rect 46147 45985 168542 46009
rect 45636 45794 164987 45818
rect 45636 45742 164849 45794
rect 164901 45742 164987 45794
rect 45636 45718 164987 45742
rect 45216 45504 161464 45528
rect 45216 45452 161304 45504
rect 161356 45452 161464 45504
rect 45216 45428 161464 45452
rect 44840 45328 157920 45352
rect 44840 45276 157763 45328
rect 157815 45276 157920 45328
rect 44840 45252 157920 45276
rect 44443 44976 154366 45000
rect 44443 44924 154216 44976
rect 154268 44924 154366 44976
rect 44443 44900 154366 44924
rect 43972 44693 150817 44717
rect 43972 44641 150665 44693
rect 150717 44641 150817 44693
rect 43972 44617 150817 44641
rect 43367 44470 147263 44494
rect 43367 44418 147097 44470
rect 147149 44418 147263 44470
rect 43367 44394 147263 44418
rect 42626 44225 143739 44249
rect 42626 44173 143572 44225
rect 143624 44173 143739 44225
rect 42626 44149 143739 44173
rect 140024 43878 140124 43879
rect 42172 43855 140197 43878
rect 42172 43803 140048 43855
rect 140100 43803 140197 43855
rect 42172 43778 140197 43803
rect 41559 43622 136634 43646
rect 41559 43570 136480 43622
rect 136532 43570 136634 43622
rect 41559 43546 136634 43570
rect 41051 43380 133086 43404
rect 41051 43328 132931 43380
rect 132983 43328 133086 43380
rect 41051 43304 133086 43328
rect 40584 43162 129567 43186
rect 40584 43110 129389 43162
rect 129441 43110 129567 43162
rect 40584 43086 129567 43110
rect 40073 42860 125996 42884
rect 40073 42808 125856 42860
rect 125908 42808 125996 42860
rect 40073 42784 125996 42808
<< via1 >>
rect 95451 687770 95823 687795
rect 95451 687448 95476 687770
rect 95476 687448 95798 687770
rect 95798 687448 95823 687770
rect 95451 687423 95823 687448
rect 172234 687993 172606 688018
rect 172234 687671 172259 687993
rect 172259 687671 172581 687993
rect 172581 687671 172606 687993
rect 172234 687646 172606 687671
rect 120776 687584 121148 687609
rect 120776 687262 120801 687584
rect 120801 687262 121123 687584
rect 121123 687262 121148 687584
rect 120776 687237 121148 687262
rect 146433 687462 146805 687487
rect 146433 687140 146458 687462
rect 146458 687140 146780 687462
rect 146780 687140 146805 687462
rect 146433 687115 146805 687140
rect 216372 687553 216744 687578
rect 216372 687231 216397 687553
rect 216397 687231 216719 687553
rect 216719 687231 216744 687553
rect 216372 687206 216744 687231
rect 223353 687628 223725 687653
rect 223353 687306 223378 687628
rect 223378 687306 223700 687628
rect 223700 687306 223725 687628
rect 223353 687281 223725 687306
rect 249023 687531 249395 687556
rect 249023 687209 249048 687531
rect 249048 687209 249370 687531
rect 249370 687209 249395 687531
rect 249023 687184 249395 687209
rect 274692 687547 275064 687572
rect 274692 687225 274717 687547
rect 274717 687225 275039 687547
rect 275039 687225 275064 687547
rect 274692 687200 275064 687225
rect 300317 687583 300689 687608
rect 300317 687261 300342 687583
rect 300342 687261 300664 687583
rect 300664 687261 300689 687583
rect 300317 687236 300689 687261
rect 325953 687548 326325 687573
rect 325953 687226 325978 687548
rect 325978 687226 326300 687548
rect 326300 687226 326325 687548
rect 325953 687201 326325 687226
rect 351618 687530 351990 687555
rect 351618 687208 351643 687530
rect 351643 687208 351965 687530
rect 351965 687208 351990 687530
rect 351618 687183 351990 687208
rect 377279 687492 377651 687517
rect 377279 687170 377304 687492
rect 377304 687170 377626 687492
rect 377626 687170 377651 687492
rect 377279 687145 377651 687170
rect 412455 687609 412827 687634
rect 412455 687287 412480 687609
rect 412480 687287 412802 687609
rect 412802 687287 412827 687609
rect 412455 687262 412827 687287
rect 428581 687599 428953 687624
rect 428581 687277 428606 687599
rect 428606 687277 428928 687599
rect 428928 687277 428953 687599
rect 428581 687252 428953 687277
rect 454215 687668 454587 687693
rect 454215 687346 454240 687668
rect 454240 687346 454562 687668
rect 454562 687346 454587 687668
rect 454215 687321 454587 687346
rect 479864 687674 480236 687699
rect 479864 687352 479889 687674
rect 479889 687352 480211 687674
rect 480211 687352 480236 687674
rect 479864 687327 480236 687352
rect 189836 660429 190208 660801
rect 569028 601724 569208 601904
rect 197193 550084 197373 550264
rect 200949 550084 201129 550264
rect 200944 548809 201124 548989
rect 193941 548353 194121 548533
rect 199445 548198 199753 548378
rect 198062 539721 198242 539901
rect 201881 539213 202061 539393
rect 565481 600723 565661 600903
rect 208759 539719 208939 539899
rect 561939 599468 562119 599648
rect 417834 577585 418014 577765
rect 558400 577586 558580 577766
rect 417838 576996 418018 577176
rect 554850 576996 555030 577176
rect 417861 576269 418041 576449
rect 551301 576269 551481 576449
rect 396874 550045 397054 550225
rect 404138 550201 404318 550381
rect 407892 550202 408072 550382
rect 406512 548254 406692 548434
rect 209982 539213 210162 539393
rect 405237 539831 405417 540011
rect 408870 539379 409050 539559
rect 206384 530732 206564 530912
rect 422060 530733 422240 530913
rect 300909 525439 301089 525619
rect 480472 520610 480652 520790
rect 275097 519234 275533 519734
rect 326559 518045 326739 518225
rect 352209 510617 352389 510797
rect 454809 510416 454989 510596
rect 377867 503193 378047 503373
rect 429162 503031 429342 503211
rect 407267 494230 407447 494410
rect 95999 445951 96179 446131
rect 76134 437865 76314 438045
rect 79782 437785 79962 437786
rect 79782 437607 79819 437785
rect 79819 437607 79925 437785
rect 79925 437607 79962 437785
rect 79782 437606 79962 437607
rect 88336 435844 88516 435845
rect 88336 435666 88373 435844
rect 88373 435666 88479 435844
rect 88479 435666 88516 435844
rect 88336 435665 88516 435666
rect 80269 435645 80449 435646
rect 80269 435467 80306 435645
rect 80306 435467 80412 435645
rect 80412 435467 80449 435645
rect 80269 435466 80449 435467
rect 76151 435109 76331 435289
rect 77082 433953 77262 434133
rect 79013 433005 79193 433185
rect 76616 431180 76988 431181
rect 76616 431002 76641 431180
rect 76641 431002 76963 431180
rect 76963 431002 76988 431180
rect 76616 431001 76988 431002
rect 77414 430118 77786 430119
rect 77414 429940 77439 430118
rect 77439 429940 77761 430118
rect 77761 429940 77786 430118
rect 77414 429939 77786 429940
rect 78423 428804 78795 428805
rect 78423 428626 78448 428804
rect 78448 428626 78770 428804
rect 78770 428626 78795 428804
rect 78423 428625 78795 428626
rect 79450 427357 79822 427358
rect 79450 427179 79475 427357
rect 79475 427179 79797 427357
rect 79797 427179 79822 427357
rect 79450 427178 79822 427179
rect 76161 424525 76341 424705
rect 76176 421759 76356 421939
rect 77115 420601 77295 420781
rect 79004 419658 79184 419838
rect 76615 417837 76987 417838
rect 76615 417659 76640 417837
rect 76640 417659 76962 417837
rect 76962 417659 76987 417837
rect 76615 417658 76987 417659
rect 77414 416772 77786 416773
rect 77414 416594 77439 416772
rect 77439 416594 77761 416772
rect 77761 416594 77786 416772
rect 77414 416593 77786 416594
rect 78425 415452 78797 415453
rect 78425 415274 78450 415452
rect 78450 415274 78772 415452
rect 78772 415274 78797 415452
rect 78425 415273 78797 415274
rect 79449 414008 79821 414009
rect 79449 413830 79474 414008
rect 79474 413830 79796 414008
rect 79796 413830 79821 414008
rect 79449 413829 79821 413830
rect 76145 411181 76325 411361
rect 76176 408414 76356 408594
rect 77103 407261 77283 407441
rect 78988 406313 79168 406493
rect 76616 404492 76988 404493
rect 76616 404314 76641 404492
rect 76641 404314 76963 404492
rect 76963 404314 76988 404492
rect 76616 404313 76988 404314
rect 77414 403428 77786 403429
rect 77414 403250 77439 403428
rect 77439 403250 77761 403428
rect 77761 403250 77786 403428
rect 77414 403249 77786 403250
rect 78423 402116 78795 402117
rect 78423 401938 78448 402116
rect 78448 401938 78770 402116
rect 78770 401938 78795 402116
rect 78423 401937 78795 401938
rect 79449 400669 79821 400670
rect 79449 400491 79474 400669
rect 79474 400491 79796 400669
rect 79796 400491 79821 400669
rect 79449 400490 79821 400491
rect 76158 397826 76338 398006
rect 76163 395072 76343 395252
rect 77115 393912 77295 394092
rect 79013 392973 79193 393153
rect 76616 391147 76988 391148
rect 76616 390969 76641 391147
rect 76641 390969 76963 391147
rect 76963 390969 76988 391147
rect 76616 390968 76988 390969
rect 77414 390081 77786 390082
rect 77414 389903 77439 390081
rect 77439 389903 77761 390081
rect 77761 389903 77786 390081
rect 77414 389902 77786 389903
rect 78423 388776 78795 388777
rect 78423 388598 78448 388776
rect 78448 388598 78770 388776
rect 78770 388598 78795 388776
rect 78423 388597 78795 388598
rect 79444 387320 79816 387321
rect 79444 387142 79469 387320
rect 79469 387142 79791 387320
rect 79791 387142 79816 387320
rect 79444 387141 79816 387142
rect 76133 384486 76313 384666
rect 76138 381724 76318 381904
rect 77103 380568 77283 380748
rect 78979 379626 79159 379806
rect 76616 377801 76988 377802
rect 76616 377623 76641 377801
rect 76641 377623 76963 377801
rect 76963 377623 76988 377801
rect 76616 377622 76988 377623
rect 77414 376737 77786 376738
rect 77414 376559 77439 376737
rect 77439 376559 77761 376737
rect 77761 376559 77786 376737
rect 77414 376558 77786 376559
rect 78423 375428 78795 375429
rect 78423 375250 78448 375428
rect 78448 375250 78770 375428
rect 78770 375250 78795 375428
rect 78423 375249 78795 375250
rect 79448 373973 79820 373974
rect 79448 373795 79473 373973
rect 79473 373795 79795 373973
rect 79795 373795 79820 373973
rect 79448 373794 79820 373795
rect 76153 371144 76333 371324
rect 76156 368383 76336 368563
rect 77065 367223 77245 367403
rect 78998 366277 79178 366457
rect 76615 364454 76987 364455
rect 76615 364276 76640 364454
rect 76640 364276 76962 364454
rect 76962 364276 76987 364454
rect 76615 364275 76987 364276
rect 77414 363395 77786 363396
rect 77414 363217 77439 363395
rect 77439 363217 77761 363395
rect 77761 363217 77786 363395
rect 77414 363216 77786 363217
rect 78420 362082 78792 362083
rect 78420 361904 78445 362082
rect 78445 361904 78767 362082
rect 78767 361904 78792 362082
rect 78420 361903 78792 361904
rect 79450 360635 79822 360636
rect 79450 360457 79475 360635
rect 79475 360457 79797 360635
rect 79797 360457 79822 360635
rect 79450 360456 79822 360457
rect 76143 357795 76323 357975
rect 76163 355038 76343 355218
rect 77155 353879 77335 354059
rect 79002 352937 79182 353117
rect 76615 351109 76987 351110
rect 76615 350931 76640 351109
rect 76640 350931 76962 351109
rect 76962 350931 76987 351109
rect 76615 350930 76987 350931
rect 77414 350049 77786 350050
rect 77414 349871 77439 350049
rect 77439 349871 77761 350049
rect 77761 349871 77786 350049
rect 77414 349870 77786 349871
rect 78423 348735 78795 348736
rect 78423 348557 78448 348735
rect 78448 348557 78770 348735
rect 78770 348557 78795 348735
rect 78423 348556 78795 348557
rect 79449 347286 79821 347287
rect 79449 347108 79474 347286
rect 79474 347108 79796 347286
rect 79796 347108 79821 347286
rect 79449 347107 79821 347108
rect 76110 344450 76290 344630
rect 76133 341688 76313 341868
rect 77121 340537 77301 340717
rect 79009 339588 79189 339768
rect 76615 337769 76987 337770
rect 76615 337591 76640 337769
rect 76640 337591 76962 337769
rect 76962 337591 76987 337769
rect 76615 337590 76987 337591
rect 77414 336702 77786 336703
rect 77414 336524 77439 336702
rect 77439 336524 77761 336702
rect 77761 336524 77786 336702
rect 77414 336523 77786 336524
rect 78418 335392 78790 335393
rect 78418 335214 78443 335392
rect 78443 335214 78765 335392
rect 78765 335214 78790 335392
rect 78418 335213 78790 335214
rect 79449 333943 79821 333944
rect 79449 333765 79474 333943
rect 79474 333765 79796 333943
rect 79796 333765 79821 333943
rect 79449 333764 79821 333765
rect 76153 331106 76333 331286
rect 76157 328348 76337 328528
rect 77109 327194 77289 327374
rect 79021 326240 79201 326420
rect 76616 324422 76988 324423
rect 76616 324244 76641 324422
rect 76641 324244 76963 324422
rect 76963 324244 76988 324422
rect 76616 324243 76988 324244
rect 77414 323358 77786 323359
rect 77414 323180 77439 323358
rect 77439 323180 77761 323358
rect 77761 323180 77786 323358
rect 77414 323179 77786 323180
rect 78423 322047 78795 322048
rect 78423 321869 78448 322047
rect 78448 321869 78770 322047
rect 78770 321869 78795 322047
rect 78423 321868 78795 321869
rect 79452 320595 79824 320596
rect 79452 320417 79477 320595
rect 79477 320417 79799 320595
rect 79799 320417 79824 320595
rect 79452 320416 79824 320417
rect 76165 317754 76345 317934
rect 76153 315003 76333 315183
rect 77114 313848 77294 314028
rect 78980 312902 79160 313082
rect 76614 311078 76986 311079
rect 76614 310900 76639 311078
rect 76639 310900 76961 311078
rect 76961 310900 76986 311078
rect 76614 310899 76986 310900
rect 77414 310013 77786 310014
rect 77414 309835 77439 310013
rect 77439 309835 77761 310013
rect 77761 309835 77786 310013
rect 77414 309834 77786 309835
rect 78424 308702 78796 308703
rect 78424 308524 78449 308702
rect 78449 308524 78771 308702
rect 78771 308524 78796 308702
rect 78424 308523 78796 308524
rect 79445 307250 79817 307251
rect 79445 307072 79470 307250
rect 79470 307072 79792 307250
rect 79792 307072 79817 307250
rect 79445 307071 79817 307072
rect 76148 304413 76328 304593
rect 76163 301656 76343 301836
rect 77120 300497 77300 300677
rect 78993 299551 79173 299731
rect 76616 297731 76988 297732
rect 76616 297553 76641 297731
rect 76641 297553 76963 297731
rect 76963 297553 76988 297731
rect 76616 297552 76988 297553
rect 77414 296665 77786 296666
rect 77414 296487 77439 296665
rect 77439 296487 77761 296665
rect 77761 296487 77786 296665
rect 77414 296486 77786 296487
rect 78425 295357 78797 295358
rect 78425 295179 78450 295357
rect 78450 295179 78772 295357
rect 78772 295179 78797 295357
rect 78425 295178 78797 295179
rect 79451 293905 79823 293906
rect 79451 293727 79476 293905
rect 79476 293727 79798 293905
rect 79798 293727 79823 293905
rect 79451 293726 79823 293727
rect 76148 291073 76328 291253
rect 76138 288320 76318 288500
rect 77117 287154 77297 287334
rect 78991 286208 79171 286388
rect 76616 284385 76988 284386
rect 76616 284207 76641 284385
rect 76641 284207 76963 284385
rect 76963 284207 76988 284385
rect 76616 284206 76988 284207
rect 77414 283323 77786 283324
rect 77414 283145 77439 283323
rect 77439 283145 77761 283323
rect 77761 283145 77786 283323
rect 77414 283144 77786 283145
rect 78423 282012 78795 282013
rect 78423 281834 78448 282012
rect 78448 281834 78770 282012
rect 78770 281834 78795 282012
rect 78423 281833 78795 281834
rect 79447 280567 79819 280568
rect 79447 280389 79472 280567
rect 79472 280389 79794 280567
rect 79794 280389 79819 280567
rect 79447 280388 79819 280389
rect 76156 277739 76336 277919
rect 76156 274961 76336 275141
rect 77128 273810 77308 273990
rect 78998 272869 79178 273049
rect 76615 271041 76987 271042
rect 76615 270863 76640 271041
rect 76640 270863 76962 271041
rect 76962 270863 76987 271041
rect 76615 270862 76987 270863
rect 77414 269976 77786 269977
rect 77414 269798 77439 269976
rect 77439 269798 77761 269976
rect 77761 269798 77786 269976
rect 77414 269797 77786 269798
rect 78424 268672 78796 268673
rect 78424 268494 78449 268672
rect 78449 268494 78771 268672
rect 78771 268494 78796 268672
rect 78424 268493 78796 268494
rect 79450 267214 79822 267215
rect 79450 267036 79475 267214
rect 79475 267036 79797 267214
rect 79797 267036 79822 267214
rect 79450 267035 79822 267036
rect 76167 264382 76347 264562
rect 76179 261623 76359 261803
rect 77130 260465 77310 260645
rect 78985 259518 79165 259698
rect 76615 257697 76987 257698
rect 76615 257519 76640 257697
rect 76640 257519 76962 257697
rect 76962 257519 76987 257697
rect 76615 257518 76987 257519
rect 77414 256633 77786 256634
rect 77414 256455 77439 256633
rect 77439 256455 77761 256633
rect 77761 256455 77786 256633
rect 77414 256454 77786 256455
rect 78423 255322 78795 255323
rect 78423 255144 78448 255322
rect 78448 255144 78770 255322
rect 78770 255144 78795 255322
rect 78423 255143 78795 255144
rect 121317 254610 121497 254790
rect 79450 253875 79822 253876
rect 79450 253697 79475 253875
rect 79475 253697 79797 253875
rect 79797 253697 79822 253875
rect 79450 253696 79822 253697
rect 76164 251033 76344 251213
rect 76162 248274 76342 248454
rect 77108 247118 77288 247298
rect 78999 246172 79179 246352
rect 76616 244351 76988 244352
rect 76616 244173 76641 244351
rect 76641 244173 76963 244351
rect 76963 244173 76988 244351
rect 76616 244172 76988 244173
rect 77414 243288 77786 243289
rect 77414 243110 77439 243288
rect 77439 243110 77761 243288
rect 77761 243110 77786 243288
rect 77414 243109 77786 243110
rect 78425 241972 78797 241973
rect 78425 241794 78450 241972
rect 78450 241794 78772 241972
rect 78772 241794 78797 241972
rect 78425 241793 78797 241794
rect 79451 240527 79823 240528
rect 79451 240349 79476 240527
rect 79476 240349 79798 240527
rect 79798 240349 79823 240527
rect 79451 240348 79823 240349
rect 76211 237660 76391 237840
rect 76209 234892 76389 235072
rect 77086 233736 77266 233916
rect 78994 232790 79174 232970
rect 76617 230968 76989 230969
rect 76617 230790 76642 230968
rect 76642 230790 76964 230968
rect 76964 230790 76989 230968
rect 76617 230789 76989 230790
rect 77414 229909 77786 229910
rect 77414 229731 77439 229909
rect 77439 229731 77761 229909
rect 77761 229731 77786 229909
rect 77414 229730 77786 229731
rect 78421 228598 78793 228599
rect 78421 228420 78446 228598
rect 78446 228420 78768 228598
rect 78768 228420 78793 228598
rect 78421 228419 78793 228420
rect 79445 227146 79817 227147
rect 79445 226968 79470 227146
rect 79470 226968 79792 227146
rect 79792 226968 79817 227146
rect 79445 226967 79817 226968
rect 93801 216514 93981 216539
rect 93801 216192 93838 216514
rect 93838 216192 93944 216514
rect 93944 216192 93981 216514
rect 93801 216167 93981 216192
rect 106151 216513 106331 216538
rect 106151 216191 106188 216513
rect 106188 216191 106294 216513
rect 106294 216191 106331 216513
rect 106151 216166 106331 216191
rect 119112 216515 119292 216540
rect 119112 216193 119149 216515
rect 119149 216193 119255 216515
rect 119255 216193 119292 216515
rect 119112 216168 119292 216193
rect 131456 216513 131636 216538
rect 131456 216191 131493 216513
rect 131493 216191 131599 216513
rect 131599 216191 131636 216513
rect 131456 216166 131636 216191
rect 144763 216512 144943 216537
rect 144763 216190 144800 216512
rect 144800 216190 144906 216512
rect 144906 216190 144943 216512
rect 144763 216165 144943 216190
rect 157106 216513 157286 216538
rect 157106 216191 157143 216513
rect 157143 216191 157249 216513
rect 157249 216191 157286 216513
rect 157106 216166 157286 216191
rect 170408 216513 170588 216538
rect 170408 216191 170445 216513
rect 170445 216191 170551 216513
rect 170551 216191 170588 216513
rect 170408 216166 170588 216191
rect 182755 216514 182935 216539
rect 182755 216192 182792 216514
rect 182792 216192 182898 216514
rect 182898 216192 182935 216514
rect 182755 216167 182935 216192
rect 196063 216515 196243 216540
rect 196063 216193 196100 216515
rect 196100 216193 196206 216515
rect 196206 216193 196243 216515
rect 196063 216168 196243 216193
rect 208407 216516 208587 216541
rect 208407 216194 208444 216516
rect 208444 216194 208550 216516
rect 208550 216194 208587 216516
rect 208407 216169 208587 216194
rect 221711 216518 221891 216543
rect 221711 216196 221748 216518
rect 221748 216196 221854 216518
rect 221854 216196 221891 216518
rect 221711 216171 221891 216196
rect 234062 216516 234242 216541
rect 234062 216194 234099 216516
rect 234099 216194 234205 216516
rect 234205 216194 234242 216516
rect 234062 216169 234242 216194
rect 247363 216515 247543 216540
rect 247363 216193 247400 216515
rect 247400 216193 247506 216515
rect 247506 216193 247543 216515
rect 247363 216168 247543 216193
rect 259712 216516 259892 216541
rect 259712 216194 259749 216516
rect 259749 216194 259855 216516
rect 259855 216194 259892 216516
rect 259712 216169 259892 216194
rect 273011 216509 273191 216534
rect 273011 216187 273048 216509
rect 273048 216187 273154 216509
rect 273154 216187 273191 216509
rect 273011 216162 273191 216187
rect 285357 216514 285537 216539
rect 285357 216192 285394 216514
rect 285394 216192 285500 216514
rect 285500 216192 285537 216514
rect 285357 216167 285537 216192
rect 298660 216516 298840 216541
rect 298660 216194 298697 216516
rect 298697 216194 298803 216516
rect 298803 216194 298840 216516
rect 298660 216169 298840 216194
rect 311007 216518 311187 216543
rect 311007 216196 311044 216518
rect 311044 216196 311150 216518
rect 311150 216196 311187 216518
rect 311007 216171 311187 216196
rect 324312 216509 324492 216534
rect 324312 216187 324349 216509
rect 324349 216187 324455 216509
rect 324455 216187 324492 216509
rect 324312 216162 324492 216187
rect 336657 216515 336837 216540
rect 336657 216193 336694 216515
rect 336694 216193 336800 216515
rect 336800 216193 336837 216515
rect 336657 216168 336837 216193
rect 349963 216513 350143 216538
rect 349963 216191 350000 216513
rect 350000 216191 350106 216513
rect 350106 216191 350143 216513
rect 349963 216166 350143 216191
rect 362308 216517 362488 216542
rect 362308 216195 362345 216517
rect 362345 216195 362451 216517
rect 362451 216195 362488 216517
rect 362308 216170 362488 216195
rect 375606 216509 375786 216534
rect 375606 216187 375643 216509
rect 375643 216187 375749 216509
rect 375749 216187 375786 216509
rect 375606 216162 375786 216187
rect 387955 216509 388135 216534
rect 387955 216187 387992 216509
rect 387992 216187 388098 216509
rect 388098 216187 388135 216509
rect 387955 216162 388135 216187
rect 401262 216512 401442 216537
rect 401262 216190 401299 216512
rect 401299 216190 401405 216512
rect 401405 216190 401442 216512
rect 401262 216165 401442 216190
rect 413612 216513 413792 216538
rect 413612 216191 413649 216513
rect 413649 216191 413755 216513
rect 413755 216191 413792 216513
rect 413612 216166 413792 216191
rect 426912 216514 427092 216539
rect 426912 216192 426949 216514
rect 426949 216192 427055 216514
rect 427055 216192 427092 216514
rect 426912 216167 427092 216192
rect 439256 216515 439436 216540
rect 439256 216193 439293 216515
rect 439293 216193 439399 216515
rect 439399 216193 439436 216515
rect 439256 216168 439436 216193
rect 452566 216524 452746 216549
rect 452566 216202 452603 216524
rect 452603 216202 452709 216524
rect 452709 216202 452746 216524
rect 452566 216177 452746 216202
rect 464906 216514 465086 216539
rect 464906 216192 464943 216514
rect 464943 216192 465049 216514
rect 465049 216192 465086 216514
rect 464906 216167 465086 216192
rect 478211 216516 478391 216541
rect 478211 216194 478248 216516
rect 478248 216194 478354 216516
rect 478354 216194 478391 216516
rect 478211 216169 478391 216194
rect 490553 216510 490733 216535
rect 490553 216188 490590 216510
rect 490590 216188 490696 216510
rect 490696 216188 490733 216510
rect 490553 216163 490733 216188
rect 94858 215760 95038 215785
rect 94858 215438 94895 215760
rect 94895 215438 95001 215760
rect 95001 215438 95038 215760
rect 94858 215413 95038 215438
rect 107208 215760 107388 215785
rect 107208 215438 107245 215760
rect 107245 215438 107351 215760
rect 107351 215438 107388 215760
rect 107208 215413 107388 215438
rect 120173 215760 120353 215785
rect 120173 215438 120210 215760
rect 120210 215438 120316 215760
rect 120316 215438 120353 215760
rect 120173 215413 120353 215438
rect 132517 215757 132697 215782
rect 132517 215435 132554 215757
rect 132554 215435 132660 215757
rect 132660 215435 132697 215757
rect 132517 215410 132697 215435
rect 145824 215760 146004 215785
rect 145824 215438 145861 215760
rect 145861 215438 145967 215760
rect 145967 215438 146004 215760
rect 145824 215413 146004 215438
rect 158164 215753 158344 215778
rect 158164 215431 158201 215753
rect 158201 215431 158307 215753
rect 158307 215431 158344 215753
rect 158164 215406 158344 215431
rect 171474 215759 171654 215784
rect 171474 215437 171511 215759
rect 171511 215437 171617 215759
rect 171617 215437 171654 215759
rect 171474 215412 171654 215437
rect 183817 215760 183997 215785
rect 183817 215438 183854 215760
rect 183854 215438 183960 215760
rect 183960 215438 183997 215760
rect 183817 215413 183997 215438
rect 197120 215761 197300 215786
rect 197120 215439 197157 215761
rect 197157 215439 197263 215761
rect 197263 215439 197300 215761
rect 197120 215414 197300 215439
rect 209468 215761 209648 215786
rect 209468 215439 209505 215761
rect 209505 215439 209611 215761
rect 209611 215439 209648 215761
rect 209468 215414 209648 215439
rect 222774 215761 222954 215786
rect 222774 215439 222811 215761
rect 222811 215439 222917 215761
rect 222917 215439 222954 215761
rect 222774 215414 222954 215439
rect 235117 215761 235297 215786
rect 235117 215439 235154 215761
rect 235154 215439 235260 215761
rect 235260 215439 235297 215761
rect 235117 215414 235297 215439
rect 248419 215760 248599 215785
rect 248419 215438 248456 215760
rect 248456 215438 248562 215760
rect 248562 215438 248599 215760
rect 248419 215413 248599 215438
rect 260770 215761 260950 215786
rect 260770 215439 260807 215761
rect 260807 215439 260913 215761
rect 260913 215439 260950 215761
rect 260770 215414 260950 215439
rect 274071 215759 274251 215784
rect 274071 215437 274108 215759
rect 274108 215437 274214 215759
rect 274214 215437 274251 215759
rect 274071 215412 274251 215437
rect 286415 215759 286595 215784
rect 286415 215437 286452 215759
rect 286452 215437 286558 215759
rect 286558 215437 286595 215759
rect 286415 215412 286595 215437
rect 299719 215761 299899 215786
rect 299719 215439 299756 215761
rect 299756 215439 299862 215761
rect 299862 215439 299899 215761
rect 299719 215414 299899 215439
rect 312066 215761 312246 215786
rect 312066 215439 312103 215761
rect 312103 215439 312209 215761
rect 312209 215439 312246 215761
rect 312066 215414 312246 215439
rect 325371 215759 325551 215784
rect 325371 215437 325408 215759
rect 325408 215437 325514 215759
rect 325514 215437 325551 215759
rect 325371 215412 325551 215437
rect 337716 215756 337896 215781
rect 337716 215434 337753 215756
rect 337753 215434 337859 215756
rect 337859 215434 337896 215756
rect 337716 215409 337896 215434
rect 351018 215759 351198 215784
rect 351018 215437 351055 215759
rect 351055 215437 351161 215759
rect 351161 215437 351198 215759
rect 351018 215412 351198 215437
rect 363367 215759 363547 215784
rect 363367 215437 363404 215759
rect 363404 215437 363510 215759
rect 363510 215437 363547 215759
rect 363367 215412 363547 215437
rect 376672 215756 376852 215781
rect 376672 215434 376709 215756
rect 376709 215434 376815 215756
rect 376815 215434 376852 215756
rect 376672 215409 376852 215434
rect 389014 215762 389194 215787
rect 389014 215440 389051 215762
rect 389051 215440 389157 215762
rect 389157 215440 389194 215762
rect 389014 215415 389194 215440
rect 402321 215758 402501 215783
rect 402321 215436 402358 215758
rect 402358 215436 402464 215758
rect 402464 215436 402501 215758
rect 402321 215411 402501 215436
rect 414668 215756 414848 215781
rect 414668 215434 414705 215756
rect 414705 215434 414811 215756
rect 414811 215434 414848 215756
rect 414668 215409 414848 215434
rect 427971 215763 428151 215788
rect 427971 215441 428008 215763
rect 428008 215441 428114 215763
rect 428114 215441 428151 215763
rect 427971 215416 428151 215441
rect 440316 215757 440496 215782
rect 440316 215435 440353 215757
rect 440353 215435 440459 215757
rect 440459 215435 440496 215757
rect 440316 215410 440496 215435
rect 453622 215763 453802 215788
rect 453622 215441 453659 215763
rect 453659 215441 453765 215763
rect 453765 215441 453802 215763
rect 453622 215416 453802 215441
rect 465968 215761 466148 215786
rect 465968 215439 466005 215761
rect 466005 215439 466111 215761
rect 466111 215439 466148 215761
rect 465968 215414 466148 215439
rect 479269 215759 479449 215784
rect 479269 215437 479306 215759
rect 479306 215437 479412 215759
rect 479412 215437 479449 215759
rect 479269 215412 479449 215437
rect 491616 215759 491796 215784
rect 491616 215437 491653 215759
rect 491653 215437 491759 215759
rect 491759 215437 491796 215759
rect 491616 215412 491796 215437
rect 91800 215070 91980 215250
rect 104145 215061 104325 215241
rect 117119 215083 117299 215263
rect 129454 215021 129634 215201
rect 142769 215037 142949 215217
rect 155109 215067 155289 215247
rect 168411 215024 168591 215204
rect 180765 215055 180945 215235
rect 194054 215083 194234 215263
rect 206412 215061 206592 215241
rect 219709 215060 219889 215240
rect 232056 215095 232236 215275
rect 245360 215079 245540 215259
rect 257705 215110 257885 215290
rect 271014 215091 271194 215271
rect 283357 215073 283537 215253
rect 296660 215069 296840 215249
rect 309004 215076 309184 215256
rect 322311 215053 322491 215233
rect 334655 215083 334835 215263
rect 347961 215053 348141 215233
rect 360305 215065 360485 215245
rect 373610 215057 373790 215237
rect 385955 215084 386135 215264
rect 399260 215083 399440 215263
rect 411609 215049 411789 215229
rect 424909 215052 425089 215232
rect 437257 215070 437437 215250
rect 450553 215070 450733 215250
rect 462904 215057 463084 215237
rect 476216 215045 476396 215225
rect 488557 215063 488737 215243
rect 96175 214879 96355 214904
rect 96175 214557 96212 214879
rect 96212 214557 96318 214879
rect 96318 214557 96355 214879
rect 96175 214532 96355 214557
rect 108518 214882 108698 214907
rect 108518 214560 108555 214882
rect 108555 214560 108661 214882
rect 108661 214560 108698 214882
rect 108518 214535 108698 214560
rect 121484 214876 121664 214901
rect 121484 214554 121521 214876
rect 121521 214554 121627 214876
rect 121627 214554 121664 214876
rect 121484 214529 121664 214554
rect 133828 214878 134008 214903
rect 133828 214556 133865 214878
rect 133865 214556 133971 214878
rect 133971 214556 134008 214878
rect 133828 214531 134008 214556
rect 147132 214878 147312 214903
rect 147132 214556 147169 214878
rect 147169 214556 147275 214878
rect 147275 214556 147312 214878
rect 147132 214531 147312 214556
rect 159480 214881 159660 214906
rect 159480 214559 159517 214881
rect 159517 214559 159623 214881
rect 159623 214559 159660 214881
rect 159480 214534 159660 214559
rect 172784 214879 172964 214904
rect 172784 214557 172821 214879
rect 172821 214557 172927 214879
rect 172927 214557 172964 214879
rect 172784 214532 172964 214557
rect 185131 214879 185311 214904
rect 185131 214557 185168 214879
rect 185168 214557 185274 214879
rect 185274 214557 185311 214879
rect 185131 214532 185311 214557
rect 198432 214877 198612 214902
rect 198432 214555 198469 214877
rect 198469 214555 198575 214877
rect 198575 214555 198612 214877
rect 198432 214530 198612 214555
rect 210781 214878 210961 214903
rect 210781 214556 210818 214878
rect 210818 214556 210924 214878
rect 210924 214556 210961 214878
rect 210781 214531 210961 214556
rect 224088 214881 224268 214906
rect 224088 214559 224125 214881
rect 224125 214559 224231 214881
rect 224231 214559 224268 214881
rect 224088 214534 224268 214559
rect 236428 214879 236608 214904
rect 236428 214557 236465 214879
rect 236465 214557 236571 214879
rect 236571 214557 236608 214879
rect 236428 214532 236608 214557
rect 249732 214876 249912 214901
rect 249732 214554 249769 214876
rect 249769 214554 249875 214876
rect 249875 214554 249912 214876
rect 249732 214529 249912 214554
rect 262080 214880 262260 214905
rect 262080 214558 262117 214880
rect 262117 214558 262223 214880
rect 262223 214558 262260 214880
rect 262080 214533 262260 214558
rect 275383 214878 275563 214903
rect 275383 214556 275420 214878
rect 275420 214556 275526 214878
rect 275526 214556 275563 214878
rect 275383 214531 275563 214556
rect 287731 214878 287911 214903
rect 287731 214556 287768 214878
rect 287768 214556 287874 214878
rect 287874 214556 287911 214878
rect 287731 214531 287911 214556
rect 301040 214881 301220 214906
rect 301040 214559 301077 214881
rect 301077 214559 301183 214881
rect 301183 214559 301220 214881
rect 301040 214534 301220 214559
rect 313378 214879 313558 214904
rect 313378 214557 313415 214879
rect 313415 214557 313521 214879
rect 313521 214557 313558 214879
rect 313378 214532 313558 214557
rect 326683 214878 326863 214903
rect 326683 214556 326720 214878
rect 326720 214556 326826 214878
rect 326826 214556 326863 214878
rect 326683 214531 326863 214556
rect 339028 214879 339208 214904
rect 339028 214557 339065 214879
rect 339065 214557 339171 214879
rect 339171 214557 339208 214879
rect 339028 214532 339208 214557
rect 352334 214876 352514 214901
rect 352334 214554 352371 214876
rect 352371 214554 352477 214876
rect 352477 214554 352514 214876
rect 352334 214529 352514 214554
rect 364679 214879 364859 214904
rect 364679 214557 364716 214879
rect 364716 214557 364822 214879
rect 364822 214557 364859 214879
rect 364679 214532 364859 214557
rect 377984 214879 378164 214904
rect 377984 214557 378021 214879
rect 378021 214557 378127 214879
rect 378127 214557 378164 214879
rect 377984 214532 378164 214557
rect 390331 214877 390511 214902
rect 390331 214555 390368 214877
rect 390368 214555 390474 214877
rect 390474 214555 390511 214877
rect 390331 214530 390511 214555
rect 403624 214869 403804 214894
rect 403624 214547 403661 214869
rect 403661 214547 403767 214869
rect 403767 214547 403804 214869
rect 403624 214522 403804 214547
rect 415976 214873 416156 214898
rect 415976 214551 416013 214873
rect 416013 214551 416119 214873
rect 416119 214551 416156 214873
rect 415976 214526 416156 214551
rect 429286 214876 429466 214901
rect 429286 214554 429323 214876
rect 429323 214554 429429 214876
rect 429429 214554 429466 214876
rect 429286 214529 429466 214554
rect 441628 214879 441808 214904
rect 441628 214557 441665 214879
rect 441665 214557 441771 214879
rect 441771 214557 441808 214879
rect 441628 214532 441808 214557
rect 454934 214882 455114 214907
rect 454934 214560 454971 214882
rect 454971 214560 455077 214882
rect 455077 214560 455114 214882
rect 454934 214535 455114 214560
rect 467278 214877 467458 214902
rect 467278 214555 467315 214877
rect 467315 214555 467421 214877
rect 467421 214555 467458 214877
rect 467278 214530 467458 214555
rect 480579 214876 480759 214901
rect 480579 214554 480616 214876
rect 480616 214554 480722 214876
rect 480722 214554 480759 214876
rect 480579 214529 480759 214554
rect 492932 214877 493112 214902
rect 492932 214555 492969 214877
rect 492969 214555 493075 214877
rect 493075 214555 493112 214877
rect 492932 214530 493112 214555
rect 97623 214090 97803 214115
rect 97623 213768 97660 214090
rect 97660 213768 97766 214090
rect 97766 213768 97803 214090
rect 97623 213743 97803 213768
rect 109981 214086 110161 214111
rect 109981 213764 110018 214086
rect 110018 213764 110124 214086
rect 110124 213764 110161 214086
rect 109981 213739 110161 213764
rect 122935 214091 123115 214116
rect 122935 213769 122972 214091
rect 122972 213769 123078 214091
rect 123078 213769 123115 214091
rect 122935 213744 123115 213769
rect 135298 214088 135478 214113
rect 135298 213766 135335 214088
rect 135335 213766 135441 214088
rect 135441 213766 135478 214088
rect 135298 213741 135478 213766
rect 148591 214080 148771 214105
rect 148591 213758 148628 214080
rect 148628 213758 148734 214080
rect 148734 213758 148771 214080
rect 148591 213733 148771 213758
rect 160931 214080 161111 214105
rect 160931 213758 160968 214080
rect 160968 213758 161074 214080
rect 161074 213758 161111 214080
rect 160931 213733 161111 213758
rect 174235 214086 174415 214111
rect 174235 213764 174272 214086
rect 174272 213764 174378 214086
rect 174378 213764 174415 214086
rect 174235 213739 174415 213764
rect 186595 214098 186775 214123
rect 186595 213776 186632 214098
rect 186632 213776 186738 214098
rect 186738 213776 186775 214098
rect 186595 213751 186775 213776
rect 199887 214080 200067 214105
rect 199887 213758 199924 214080
rect 199924 213758 200030 214080
rect 200030 213758 200067 214080
rect 199887 213733 200067 213758
rect 212236 214094 212416 214119
rect 212236 213772 212273 214094
rect 212273 213772 212379 214094
rect 212379 213772 212416 214094
rect 212236 213747 212416 213772
rect 225542 214088 225722 214113
rect 225542 213766 225579 214088
rect 225579 213766 225685 214088
rect 225685 213766 225722 214088
rect 225542 213741 225722 213766
rect 237896 214090 238076 214115
rect 237896 213768 237933 214090
rect 237933 213768 238039 214090
rect 238039 213768 238076 214090
rect 237896 213743 238076 213768
rect 251199 214091 251379 214116
rect 251199 213769 251236 214091
rect 251236 213769 251342 214091
rect 251342 213769 251379 214091
rect 251199 213744 251379 213769
rect 263541 214095 263721 214120
rect 263541 213773 263578 214095
rect 263578 213773 263684 214095
rect 263684 213773 263721 214095
rect 263541 213748 263721 213773
rect 276848 214086 277028 214111
rect 276848 213764 276885 214086
rect 276885 213764 276991 214086
rect 276991 213764 277028 214086
rect 276848 213739 277028 213764
rect 289177 214085 289357 214110
rect 289177 213763 289214 214085
rect 289214 213763 289320 214085
rect 289320 213763 289357 214085
rect 289177 213738 289357 213763
rect 302496 214088 302676 214113
rect 302496 213766 302533 214088
rect 302533 213766 302639 214088
rect 302639 213766 302676 214088
rect 302496 213741 302676 213766
rect 314835 214091 315015 214116
rect 314835 213769 314872 214091
rect 314872 213769 314978 214091
rect 314978 213769 315015 214091
rect 314835 213744 315015 213769
rect 328133 214091 328313 214116
rect 328133 213769 328170 214091
rect 328170 213769 328276 214091
rect 328276 213769 328313 214091
rect 328133 213744 328313 213769
rect 340483 214092 340663 214117
rect 340483 213770 340520 214092
rect 340520 213770 340626 214092
rect 340626 213770 340663 214092
rect 340483 213745 340663 213770
rect 353792 214088 353972 214113
rect 353792 213766 353829 214088
rect 353829 213766 353935 214088
rect 353935 213766 353972 214088
rect 353792 213741 353972 213766
rect 366126 214093 366306 214118
rect 366126 213771 366163 214093
rect 366163 213771 366269 214093
rect 366269 213771 366306 214093
rect 366126 213746 366306 213771
rect 379444 214092 379624 214117
rect 379444 213770 379481 214092
rect 379481 213770 379587 214092
rect 379587 213770 379624 214092
rect 379444 213745 379624 213770
rect 391778 214089 391958 214114
rect 391778 213767 391815 214089
rect 391815 213767 391921 214089
rect 391921 213767 391958 214089
rect 391778 213742 391958 213767
rect 405089 214085 405269 214110
rect 405089 213763 405126 214085
rect 405126 213763 405232 214085
rect 405232 213763 405269 214085
rect 405089 213738 405269 213763
rect 417437 214095 417617 214120
rect 417437 213773 417474 214095
rect 417474 213773 417580 214095
rect 417580 213773 417617 214095
rect 417437 213748 417617 213773
rect 430752 214094 430932 214119
rect 430752 213772 430789 214094
rect 430789 213772 430895 214094
rect 430895 213772 430932 214094
rect 430752 213747 430932 213772
rect 443088 214088 443268 214113
rect 443088 213766 443125 214088
rect 443125 213766 443231 214088
rect 443231 213766 443268 214088
rect 443088 213741 443268 213766
rect 456393 214088 456573 214113
rect 456393 213766 456430 214088
rect 456430 213766 456536 214088
rect 456536 213766 456573 214088
rect 456393 213741 456573 213766
rect 468746 214094 468926 214119
rect 468746 213772 468783 214094
rect 468783 213772 468889 214094
rect 468889 213772 468926 214094
rect 468746 213747 468926 213772
rect 482048 214088 482228 214113
rect 482048 213766 482085 214088
rect 482085 213766 482191 214088
rect 482191 213766 482228 214088
rect 482048 213741 482228 213766
rect 494383 214089 494563 214114
rect 494383 213767 494420 214089
rect 494420 213767 494526 214089
rect 494526 213767 494563 214089
rect 494383 213742 494563 213767
rect 90853 213265 91033 213445
rect 103203 213263 103383 213443
rect 116163 213264 116343 213444
rect 128506 213223 128686 213403
rect 141811 213183 141991 213363
rect 154155 213248 154335 213428
rect 167466 213209 167646 213389
rect 179810 213243 179990 213423
rect 193120 213235 193300 213415
rect 205456 213249 205636 213429
rect 218761 213250 218941 213430
rect 231111 213237 231291 213417
rect 244410 213227 244590 213407
rect 256759 213247 256939 213427
rect 270068 213228 270248 213408
rect 282412 213205 282592 213385
rect 295715 213220 295895 213400
rect 308063 213178 308243 213358
rect 321361 213237 321541 213417
rect 333706 213194 333886 213374
rect 347012 213261 347192 213441
rect 359361 213249 359541 213429
rect 372664 213261 372844 213441
rect 385011 213262 385191 213442
rect 398308 213257 398488 213437
rect 410656 213257 410836 213437
rect 423965 213260 424145 213440
rect 436214 213157 436586 213529
rect 449615 213253 449795 213433
rect 461963 213251 462143 213431
rect 475260 213246 475440 213426
rect 487608 213220 487788 213400
rect 86939 212604 87119 212784
rect 89701 212573 89881 212753
rect 99284 212553 99464 212733
rect 102057 212578 102237 212758
rect 112244 212588 112424 212768
rect 115011 212613 115191 212793
rect 124583 212578 124763 212758
rect 127356 212569 127536 212749
rect 137899 212565 138079 212745
rect 140661 212585 140841 212765
rect 150241 212526 150421 212706
rect 152999 212542 153179 212722
rect 163541 212543 163721 212723
rect 166312 212531 166492 212711
rect 175891 212550 176071 212730
rect 178652 212531 178832 212711
rect 189195 212557 189375 212737
rect 191962 212557 192142 212737
rect 201536 212567 201716 212747
rect 204302 212545 204482 212725
rect 214844 212587 215024 212767
rect 217608 212583 217788 212763
rect 227195 212576 227375 212756
rect 229954 212554 230134 212734
rect 240496 212575 240676 212755
rect 243257 212584 243437 212764
rect 252842 212565 253022 212745
rect 255602 212565 255782 212745
rect 266143 212481 266323 212661
rect 268910 212515 269090 212695
rect 278487 212546 278667 212726
rect 281255 212556 281435 212736
rect 291795 212490 291975 212670
rect 294558 212511 294738 212691
rect 304147 212531 304327 212711
rect 306911 212526 307091 212706
rect 317450 212546 317630 212726
rect 320208 212546 320388 212726
rect 329791 212573 329971 212753
rect 332554 212608 332734 212788
rect 343097 212544 343277 212724
rect 345859 212549 346039 212729
rect 355438 212540 355618 212720
rect 358204 212559 358384 212739
rect 368747 212526 368927 212706
rect 371509 212550 371689 212730
rect 381091 212573 381271 212753
rect 383856 212592 384036 212772
rect 394398 212537 394578 212717
rect 397159 212587 397339 212767
rect 406737 212553 406917 212733
rect 409506 212573 409686 212753
rect 420047 212578 420227 212758
rect 422810 212596 422990 212776
rect 432396 212593 432576 212773
rect 435155 212565 435335 212745
rect 445691 212510 445871 212690
rect 448459 212564 448639 212744
rect 458041 212525 458221 212705
rect 460803 212557 460983 212737
rect 471338 212479 471518 212659
rect 474110 212533 474290 212713
rect 483694 212491 483874 212671
rect 486457 212561 486637 212741
rect 292516 78843 292568 78895
rect 288955 77783 289007 77835
rect 285422 76732 285474 76784
rect 281872 75085 281924 75137
rect 278312 74267 278364 74319
rect 274773 73190 274825 73242
rect 271233 71845 271285 71897
rect 267693 70469 267745 70521
rect 264145 69582 264197 69634
rect 260593 67230 260645 67282
rect 257049 66596 257101 66648
rect 253511 65300 253563 65352
rect 249945 64146 249997 64198
rect 246384 63303 246436 63355
rect 242866 62475 242918 62527
rect 239313 61741 239365 61793
rect 179041 46789 179093 46841
rect 175484 46513 175536 46565
rect 171955 46248 172007 46300
rect 168401 46009 168453 46061
rect 164849 45742 164901 45794
rect 161304 45452 161356 45504
rect 157763 45276 157815 45328
rect 154216 44924 154268 44976
rect 150665 44641 150717 44693
rect 147097 44418 147149 44470
rect 143572 44173 143624 44225
rect 140048 43803 140100 43855
rect 136480 43570 136532 43622
rect 132931 43328 132983 43380
rect 129389 43110 129441 43162
rect 125856 42808 125908 42860
<< metal2 >>
rect 538244 694820 538644 694956
rect 538244 694684 538383 694820
rect 538519 694684 538644 694820
rect 172220 688020 172620 688032
rect 95437 687797 95837 687809
rect 95437 687421 95449 687797
rect 95825 687421 95837 687797
rect 172220 687644 172232 688020
rect 172608 687644 172620 688020
rect 454201 687695 454601 687707
rect 172220 687632 172620 687644
rect 223339 687655 223739 687667
rect 95437 687409 95837 687421
rect 120762 687611 121162 687623
rect 120762 687235 120774 687611
rect 121150 687235 121162 687611
rect 216358 687580 216758 687592
rect 120762 687223 121162 687235
rect 146419 687489 146819 687501
rect 146419 687113 146431 687489
rect 146807 687113 146819 687489
rect 216358 687204 216370 687580
rect 216746 687204 216758 687580
rect 223339 687279 223351 687655
rect 223727 687279 223739 687655
rect 412441 687636 412841 687648
rect 300303 687610 300703 687622
rect 274678 687574 275078 687586
rect 223339 687267 223739 687279
rect 249009 687558 249409 687570
rect 216358 687192 216758 687204
rect 249009 687182 249021 687558
rect 249397 687182 249409 687558
rect 274678 687198 274690 687574
rect 275066 687198 275078 687574
rect 300303 687234 300315 687610
rect 300691 687234 300703 687610
rect 300303 687222 300703 687234
rect 325939 687575 326339 687587
rect 274678 687186 275078 687198
rect 325939 687199 325951 687575
rect 326327 687199 326339 687575
rect 325939 687187 326339 687199
rect 351604 687557 352004 687569
rect 249009 687170 249409 687182
rect 351604 687181 351616 687557
rect 351992 687181 352004 687557
rect 351604 687169 352004 687181
rect 377265 687519 377665 687531
rect 377265 687143 377277 687519
rect 377653 687143 377665 687519
rect 412441 687260 412453 687636
rect 412829 687260 412841 687636
rect 412441 687248 412841 687260
rect 428567 687626 428967 687638
rect 428567 687250 428579 687626
rect 428955 687250 428967 687626
rect 454201 687319 454213 687695
rect 454589 687319 454601 687695
rect 454201 687307 454601 687319
rect 479850 687701 480250 687713
rect 479850 687325 479862 687701
rect 480238 687325 480250 687701
rect 479850 687313 480250 687325
rect 428567 687238 428967 687250
rect 377265 687131 377665 687143
rect 146419 687101 146819 687113
rect 538244 674838 538644 694684
rect 198417 674686 538644 674838
rect 198417 674550 198548 674686
rect 198684 674550 538644 674686
rect 198417 674438 538644 674550
rect 19989 660806 20389 660809
rect 189822 660806 190222 660815
rect 19905 660801 397363 660806
rect 19905 660797 189836 660801
rect 19905 660421 20001 660797
rect 20377 660429 189836 660797
rect 190208 660679 397363 660801
rect 190208 660543 396896 660679
rect 397032 660543 397363 660679
rect 190208 660429 397363 660543
rect 20377 660421 397363 660429
rect 19905 660406 397363 660421
rect 416056 659178 436197 659190
rect 416056 658802 416192 659178
rect 416568 658802 436197 659178
rect 416056 658790 436197 658802
rect 414171 577765 418162 577776
rect 414171 577585 417834 577765
rect 418014 577585 418162 577765
rect 414171 577576 418162 577585
rect 4997 560743 390842 560757
rect 4997 560367 5039 560743
rect 5415 560367 390842 560743
rect 4997 560357 390842 560367
rect 5027 560355 5427 560357
rect 181965 559703 182460 559735
rect 181965 559327 182013 559703
rect 182389 559327 182460 559703
rect 181965 559293 182460 559327
rect 183496 559311 183896 560357
rect 388949 559763 389349 559775
rect 184993 559671 185393 559683
rect 184993 559295 185005 559671
rect 185381 559295 185393 559671
rect 184993 559283 185393 559295
rect 186484 559680 186884 559692
rect 186484 559304 186496 559680
rect 186872 559304 186884 559680
rect 186484 559292 186884 559304
rect 198418 559579 198818 559591
rect 198418 559203 198430 559579
rect 198806 559203 198818 559579
rect 388949 559387 388961 559763
rect 389337 559387 389349 559763
rect 388949 559375 389349 559387
rect 390442 559366 390842 560357
rect 391996 559679 392396 559691
rect 391996 559303 392008 559679
rect 392384 559303 392396 559679
rect 391996 559291 392396 559303
rect 393428 559665 393828 559677
rect 393428 559289 393440 559665
rect 393816 559289 393828 559665
rect 393428 559277 393828 559289
rect 405352 559664 405752 559676
rect 405352 559288 405364 559664
rect 405740 559288 405752 559664
rect 405352 559276 405752 559288
rect 198418 559191 198818 559203
rect 410969 556818 411169 556850
rect 204029 556748 204229 556780
rect 204029 556612 204061 556748
rect 204197 556612 204229 556748
rect 410969 556682 411001 556818
rect 411137 556682 411169 556818
rect 410969 556650 411169 556682
rect 204029 556580 204229 556612
rect 203981 556092 204694 556292
rect 410925 556138 411796 556338
rect 24149 553635 24549 553640
rect 24149 553623 24550 553635
rect 24149 553247 24162 553623
rect 24538 553247 24550 553623
rect 24149 553235 24550 553247
rect 24149 215789 24549 553235
rect 204494 550743 204694 556092
rect 411596 553666 411796 556138
rect 410316 553466 411796 553666
rect 203370 550543 398692 550743
rect 407882 550391 408082 550392
rect 404128 550382 408083 550391
rect 404128 550381 407892 550382
rect 197184 550274 201138 550275
rect 197183 550264 201139 550274
rect 197183 550084 197193 550264
rect 197373 550084 200949 550264
rect 201129 550084 201139 550264
rect 197183 550075 201139 550084
rect 197183 550074 197383 550075
rect 200939 550074 201139 550075
rect 396864 550225 397064 550235
rect 396864 550045 396874 550225
rect 397054 550045 397064 550225
rect 404128 550201 404138 550381
rect 404318 550202 407892 550381
rect 408072 550202 408083 550382
rect 404318 550201 408083 550202
rect 404128 550191 408083 550201
rect 396864 550035 397064 550045
rect 200934 548989 201134 548999
rect 200934 548809 200944 548989
rect 201124 548809 201134 548989
rect 200934 548799 201134 548809
rect 193931 548533 194131 548543
rect 193931 548353 193941 548533
rect 194121 548353 194131 548533
rect 406486 548462 406718 548470
rect 406400 548434 406874 548462
rect 199428 548404 199770 548416
rect 193931 548343 194131 548353
rect 199252 548378 199798 548404
rect 199252 548198 199445 548378
rect 199753 548198 199798 548378
rect 406400 548254 406512 548434
rect 406692 548254 406874 548434
rect 406400 548222 406874 548254
rect 406486 548218 406718 548222
rect 199252 548170 199798 548198
rect 199428 548160 199770 548170
rect 37851 542707 38251 542719
rect 37851 542331 37863 542707
rect 38239 542623 38251 542707
rect 38239 542423 191747 542623
rect 38239 542331 38251 542423
rect 37851 542319 38251 542331
rect 184162 530891 184362 540674
rect 184162 530755 184194 530891
rect 184330 530755 184362 530891
rect 184162 530723 184362 530755
rect 197444 530892 197644 540790
rect 198052 539901 198252 539911
rect 198052 539721 198062 539901
rect 198242 539721 198252 539901
rect 198052 539711 198252 539721
rect 208749 539899 208949 539909
rect 208749 539719 208759 539899
rect 208939 539719 208949 539899
rect 208749 539709 208949 539719
rect 201871 539393 202071 539403
rect 201871 539213 201881 539393
rect 202061 539213 202071 539393
rect 201871 539203 202071 539213
rect 209972 539393 210172 539403
rect 209972 539213 209982 539393
rect 210162 539213 210172 539393
rect 209972 539203 210172 539213
rect 197444 530756 197476 530892
rect 197612 530756 197644 530892
rect 197444 530622 197644 530756
rect 206374 530912 206574 530922
rect 206374 530732 206384 530912
rect 206564 530732 206574 530912
rect 206374 530722 206574 530732
rect 391148 530892 391348 540695
rect 391148 530756 391180 530892
rect 391316 530756 391348 530892
rect 391148 530723 391348 530756
rect 404393 530891 404593 540852
rect 414171 540682 414371 577576
rect 417824 577575 418024 577576
rect 414658 577176 418160 577186
rect 414658 576996 417838 577176
rect 418018 576996 418160 577176
rect 414658 576986 418160 576996
rect 414658 547573 414858 576986
rect 414658 547437 414690 547573
rect 414826 547437 414858 547573
rect 414658 547352 414858 547437
rect 415335 576449 418191 576459
rect 415335 576269 417861 576449
rect 418041 576269 418191 576449
rect 415335 576259 418191 576269
rect 415335 547580 415535 576259
rect 435797 550038 436197 658790
rect 569018 601904 569218 601976
rect 569018 601724 569028 601904
rect 569208 601724 569218 601904
rect 565471 600903 565671 600948
rect 565471 600723 565481 600903
rect 565661 600723 565671 600903
rect 561929 599648 562129 599685
rect 561929 599468 561939 599648
rect 562119 599468 562129 599648
rect 558390 577766 558590 577817
rect 558390 577586 558400 577766
rect 558580 577586 558590 577766
rect 554840 577176 555040 577232
rect 554840 576996 554850 577176
rect 555030 576996 555040 577176
rect 551291 576449 551491 576498
rect 551291 576269 551301 576449
rect 551481 576269 551491 576449
rect 435797 549638 497071 550038
rect 415335 547444 415367 547580
rect 415503 547444 415535 547580
rect 415335 547349 415535 547444
rect 410746 540482 414371 540682
rect 405227 540011 405427 540021
rect 405227 539831 405237 540011
rect 405417 539831 405427 540011
rect 405227 539821 405427 539831
rect 408860 539559 409060 539569
rect 408860 539379 408870 539559
rect 409050 539379 409060 539559
rect 408860 539369 409060 539379
rect 404393 530755 404425 530891
rect 404561 530755 404593 530891
rect 404393 530625 404593 530755
rect 422050 530913 422250 530923
rect 422050 530733 422060 530913
rect 422240 530733 422250 530913
rect 422050 530723 422250 530733
rect 300899 525619 301099 525629
rect 300899 525439 300909 525619
rect 301089 525439 301099 525619
rect 300899 525429 301099 525439
rect 480462 520790 480662 520800
rect 480462 520610 480472 520790
rect 480652 520610 480662 520790
rect 480462 520600 480662 520610
rect 275068 519734 275562 519754
rect 275068 519606 275097 519734
rect 275068 519234 275097 519366
rect 275533 519606 275562 519734
rect 275533 519234 275562 519366
rect 275068 519214 275562 519234
rect 326549 518225 326749 518235
rect 326549 518045 326559 518225
rect 326739 518045 326749 518225
rect 326549 518035 326749 518045
rect 352199 510797 352399 510807
rect 352199 510617 352209 510797
rect 352389 510617 352399 510797
rect 352199 510607 352399 510617
rect 454799 510596 454999 510606
rect 454799 510416 454809 510596
rect 454989 510416 454999 510596
rect 454799 510406 454999 510416
rect 377857 503373 378057 503383
rect 377857 503193 377867 503373
rect 378047 503193 378057 503373
rect 377857 503183 378057 503193
rect 429152 503211 429352 503221
rect 429152 503031 429162 503211
rect 429342 503031 429352 503211
rect 429152 503021 429352 503031
rect 407257 494410 407457 494420
rect 407257 494230 407267 494410
rect 407447 494230 407457 494410
rect 407257 494220 407457 494230
rect 95989 446131 96189 446141
rect 95989 445951 95999 446131
rect 96179 445951 96189 446131
rect 95989 445941 96189 445951
rect 76124 438045 76324 438055
rect 76124 437865 76134 438045
rect 76314 437865 76324 438045
rect 76124 437855 76324 437865
rect 79772 437786 79972 437796
rect 79772 437606 79782 437786
rect 79962 437606 79972 437786
rect 79772 437596 79972 437606
rect 48822 437001 75992 437101
rect 24149 215413 24161 215789
rect 24537 215413 24549 215789
rect 24149 215399 24549 215413
rect 29663 225136 29863 225170
rect 29663 225000 29695 225136
rect 29831 225000 29863 225136
rect 29663 124938 29863 225000
rect 216 124905 29863 124938
rect 216 124769 273 124905
rect 409 124769 29863 124905
rect 216 124738 29863 124769
rect 241 124737 441 124738
rect 48822 48694 48922 437001
rect 88326 435845 88526 435855
rect 88326 435665 88336 435845
rect 88516 435665 88526 435845
rect 80259 435646 80459 435656
rect 88326 435655 88526 435665
rect 80259 435466 80269 435646
rect 80449 435466 80459 435646
rect 80259 435456 80459 435466
rect 76141 435289 76341 435299
rect 76141 435109 76151 435289
rect 76331 435109 76341 435289
rect 76141 435099 76341 435109
rect 77072 434133 77272 434143
rect 77072 433953 77082 434133
rect 77262 433953 77272 434133
rect 77072 433943 77272 433953
rect 79003 433185 79203 433195
rect 79003 433005 79013 433185
rect 79193 433005 79203 433185
rect 79003 432995 79203 433005
rect 76601 431191 77001 431198
rect 76601 431181 77002 431191
rect 76601 431001 76616 431181
rect 76988 431001 77002 431181
rect 76601 430991 77002 431001
rect 76151 424705 76351 424715
rect 76151 424525 76161 424705
rect 76341 424525 76351 424705
rect 76151 424515 76351 424525
rect 49956 423659 75981 423759
rect 49956 49896 50056 423659
rect 76166 421939 76366 421949
rect 76166 421759 76176 421939
rect 76356 421759 76366 421939
rect 76166 421749 76366 421759
rect 76601 417838 77001 430991
rect 77400 430119 77800 430133
rect 77400 429939 77414 430119
rect 77786 429939 77800 430119
rect 77105 420781 77305 420791
rect 77105 420601 77115 420781
rect 77295 420601 77305 420781
rect 77105 420591 77305 420601
rect 76601 417658 76615 417838
rect 76987 417658 77001 417838
rect 76135 411361 76335 411371
rect 76135 411181 76145 411361
rect 76325 411181 76335 411361
rect 76135 411171 76335 411181
rect 50678 410291 75943 410391
rect 50678 50968 50778 410291
rect 76166 408594 76366 408604
rect 76166 408414 76176 408594
rect 76356 408414 76366 408594
rect 76166 408404 76366 408414
rect 76601 404503 77001 417658
rect 77400 416773 77800 429939
rect 77400 416593 77414 416773
rect 77786 416593 77800 416773
rect 77093 407441 77293 407451
rect 77093 407261 77103 407441
rect 77283 407261 77293 407441
rect 77093 407251 77293 407261
rect 76601 404493 77002 404503
rect 76601 404313 76616 404493
rect 76988 404313 77002 404493
rect 76601 404303 77002 404313
rect 76148 398006 76348 398016
rect 76148 397826 76158 398006
rect 76338 397826 76348 398006
rect 76148 397816 76348 397826
rect 51598 396961 75932 397061
rect 51598 51707 51698 396961
rect 76153 395252 76353 395262
rect 76153 395072 76163 395252
rect 76343 395072 76353 395252
rect 76153 395062 76353 395072
rect 76601 391158 77001 404303
rect 77400 403429 77800 416593
rect 77400 403249 77414 403429
rect 77786 403249 77800 403429
rect 77105 394092 77305 394102
rect 77105 393912 77115 394092
rect 77295 393912 77305 394092
rect 77105 393902 77305 393912
rect 76601 391148 77002 391158
rect 76601 390968 76616 391148
rect 76988 390968 77002 391148
rect 76601 390958 77002 390968
rect 76123 384666 76323 384676
rect 76123 384486 76133 384666
rect 76313 384486 76323 384666
rect 76123 384476 76323 384486
rect 52081 383620 75947 383720
rect 52081 52470 52181 383620
rect 76128 381904 76328 381914
rect 76128 381724 76138 381904
rect 76318 381724 76328 381904
rect 76128 381714 76328 381724
rect 76601 377812 77001 390958
rect 77400 390082 77800 403249
rect 77400 389902 77414 390082
rect 77786 389902 77800 390082
rect 77093 380748 77293 380758
rect 77093 380568 77103 380748
rect 77283 380568 77293 380748
rect 77093 380558 77293 380568
rect 76601 377802 77002 377812
rect 76601 377622 76616 377802
rect 76988 377622 77002 377802
rect 76601 377612 77002 377622
rect 76143 371324 76343 371334
rect 76143 371144 76153 371324
rect 76333 371144 76343 371324
rect 76143 371134 76343 371144
rect 52556 370277 75952 370377
rect 52556 53517 52656 370277
rect 76146 368563 76346 368573
rect 76146 368383 76156 368563
rect 76336 368383 76346 368563
rect 76146 368373 76346 368383
rect 76601 364455 77001 377612
rect 77400 376738 77800 389902
rect 77400 376558 77414 376738
rect 77786 376558 77800 376738
rect 77055 367403 77255 367413
rect 77055 367223 77065 367403
rect 77245 367223 77255 367403
rect 77055 367213 77255 367223
rect 76601 364275 76615 364455
rect 76987 364275 77001 364455
rect 76133 357975 76333 357985
rect 76133 357795 76143 357975
rect 76323 357795 76333 357975
rect 76133 357785 76333 357795
rect 52854 356944 75945 357044
rect 52854 53982 52954 356944
rect 76153 355218 76353 355228
rect 76153 355038 76163 355218
rect 76343 355038 76353 355218
rect 76153 355028 76353 355038
rect 76601 351110 77001 364275
rect 77400 363396 77800 376558
rect 77400 363216 77414 363396
rect 77786 363216 77800 363396
rect 77145 354059 77345 354069
rect 77145 353879 77155 354059
rect 77335 353879 77345 354059
rect 77145 353869 77345 353879
rect 76601 350930 76615 351110
rect 76987 350930 77001 351110
rect 76100 344630 76300 344640
rect 76100 344450 76110 344630
rect 76290 344450 76300 344630
rect 76100 344440 76300 344450
rect 53197 343591 75937 343691
rect 53197 54695 53297 343591
rect 76123 341868 76323 341878
rect 76123 341688 76133 341868
rect 76313 341688 76323 341868
rect 76123 341678 76323 341688
rect 76601 337770 77001 350930
rect 77400 350050 77800 363216
rect 78409 428805 78809 428821
rect 78409 428625 78423 428805
rect 78795 428625 78809 428805
rect 78409 415463 78809 428625
rect 79433 427368 79833 427384
rect 79433 427358 79836 427368
rect 79433 427178 79450 427358
rect 79822 427178 79836 427358
rect 79433 427168 79836 427178
rect 78994 419838 79194 419848
rect 78994 419658 79004 419838
rect 79184 419658 79194 419838
rect 78994 419648 79194 419658
rect 78409 415453 78811 415463
rect 78409 415273 78425 415453
rect 78797 415273 78811 415453
rect 78409 415263 78811 415273
rect 78409 402117 78809 415263
rect 79433 414019 79833 427168
rect 79433 414009 79835 414019
rect 79433 413829 79449 414009
rect 79821 413829 79835 414009
rect 79433 413819 79835 413829
rect 78978 406493 79178 406503
rect 78978 406313 78988 406493
rect 79168 406313 79178 406493
rect 78978 406303 79178 406313
rect 78409 401937 78423 402117
rect 78795 401937 78809 402117
rect 78409 388777 78809 401937
rect 79433 400680 79833 413819
rect 79433 400670 79835 400680
rect 79433 400490 79449 400670
rect 79821 400490 79835 400670
rect 79433 400480 79835 400490
rect 79003 393153 79203 393163
rect 79003 392973 79013 393153
rect 79193 392973 79203 393153
rect 79003 392963 79203 392973
rect 78409 388597 78423 388777
rect 78795 388597 78809 388777
rect 78409 375429 78809 388597
rect 79433 387331 79833 400480
rect 79430 387321 79833 387331
rect 79430 387141 79444 387321
rect 79816 387141 79833 387321
rect 79430 387131 79833 387141
rect 78969 379806 79169 379816
rect 78969 379626 78979 379806
rect 79159 379626 79169 379806
rect 78969 379616 79169 379626
rect 78409 375249 78423 375429
rect 78795 375249 78809 375429
rect 78409 362093 78809 375249
rect 79433 373984 79833 387131
rect 79433 373974 79834 373984
rect 79433 373794 79448 373974
rect 79820 373794 79834 373974
rect 79433 373784 79834 373794
rect 78988 366457 79188 366467
rect 78988 366277 78998 366457
rect 79178 366277 79188 366457
rect 78988 366267 79188 366277
rect 78406 362083 78809 362093
rect 78406 361903 78420 362083
rect 78792 361903 78809 362083
rect 78406 361893 78809 361903
rect 77400 349870 77414 350050
rect 77786 349870 77800 350050
rect 77111 340717 77311 340727
rect 77111 340537 77121 340717
rect 77301 340537 77311 340717
rect 77111 340527 77311 340537
rect 76601 337590 76615 337770
rect 76987 337590 77001 337770
rect 76143 331286 76343 331296
rect 76143 331106 76153 331286
rect 76333 331106 76343 331286
rect 76143 331096 76343 331106
rect 53572 330245 75955 330345
rect 53572 55175 53672 330245
rect 76147 328528 76347 328538
rect 76147 328348 76157 328528
rect 76337 328348 76347 328528
rect 76147 328338 76347 328348
rect 76601 324433 77001 337590
rect 77400 336703 77800 349870
rect 77400 336523 77414 336703
rect 77786 336523 77800 336703
rect 77099 327374 77299 327384
rect 77099 327194 77109 327374
rect 77289 327194 77299 327374
rect 77099 327184 77299 327194
rect 76601 324423 77002 324433
rect 76601 324243 76616 324423
rect 76988 324243 77002 324423
rect 76601 324233 77002 324243
rect 76155 317934 76355 317944
rect 76155 317754 76165 317934
rect 76345 317754 76355 317934
rect 76155 317744 76355 317754
rect 53978 316895 75959 316995
rect 53978 55699 54078 316895
rect 76143 315183 76343 315193
rect 76143 315003 76153 315183
rect 76333 315003 76343 315183
rect 76143 314993 76343 315003
rect 76601 311089 77001 324233
rect 77400 323359 77800 336523
rect 78409 348736 78809 361893
rect 79433 360646 79833 373784
rect 79433 360636 79836 360646
rect 79433 360456 79450 360636
rect 79822 360456 79836 360636
rect 79433 360446 79836 360456
rect 78992 353117 79192 353127
rect 78992 352937 79002 353117
rect 79182 352937 79192 353117
rect 78992 352927 79192 352937
rect 78409 348556 78423 348736
rect 78795 348556 78809 348736
rect 78409 335403 78809 348556
rect 79433 347297 79833 360446
rect 79433 347287 79835 347297
rect 79433 347107 79449 347287
rect 79821 347107 79835 347287
rect 79433 347097 79835 347107
rect 78999 339768 79199 339778
rect 78999 339588 79009 339768
rect 79189 339588 79199 339768
rect 78999 339578 79199 339588
rect 78404 335393 78809 335403
rect 78404 335213 78418 335393
rect 78790 335213 78809 335393
rect 78404 335203 78809 335213
rect 77400 323179 77414 323359
rect 77786 323179 77800 323359
rect 77104 314028 77304 314038
rect 77104 313848 77114 314028
rect 77294 313848 77304 314028
rect 77104 313838 77304 313848
rect 76600 311079 77001 311089
rect 76600 310899 76614 311079
rect 76986 310899 77001 311079
rect 76600 310889 77001 310899
rect 76138 304593 76338 304603
rect 76138 304413 76148 304593
rect 76328 304413 76338 304593
rect 76138 304403 76338 304413
rect 54315 303544 75942 303644
rect 54315 56057 54415 303544
rect 76153 301836 76353 301846
rect 76153 301656 76163 301836
rect 76343 301656 76353 301836
rect 76153 301646 76353 301656
rect 76601 297742 77001 310889
rect 77400 310014 77800 323179
rect 77400 309834 77414 310014
rect 77786 309834 77800 310014
rect 77110 300677 77310 300687
rect 77110 300497 77120 300677
rect 77300 300497 77310 300677
rect 77110 300487 77310 300497
rect 76601 297732 77002 297742
rect 76601 297552 76616 297732
rect 76988 297552 77002 297732
rect 76601 297542 77002 297552
rect 76138 291253 76338 291263
rect 76138 291073 76148 291253
rect 76328 291073 76338 291253
rect 76138 291063 76338 291073
rect 54700 290206 75952 290306
rect 54700 56341 54800 290206
rect 76128 288500 76328 288510
rect 76128 288320 76138 288500
rect 76318 288320 76328 288500
rect 76128 288310 76328 288320
rect 76601 284396 77001 297542
rect 77400 296666 77800 309834
rect 77400 296486 77414 296666
rect 77786 296486 77800 296666
rect 77107 287334 77307 287344
rect 77107 287154 77117 287334
rect 77297 287154 77307 287334
rect 77107 287144 77307 287154
rect 76601 284386 77002 284396
rect 76601 284206 76616 284386
rect 76988 284206 77002 284386
rect 76601 284196 77002 284206
rect 76146 277919 76346 277929
rect 76146 277739 76156 277919
rect 76336 277739 76346 277919
rect 76146 277729 76346 277739
rect 54958 276865 75939 276965
rect 54958 56748 55058 276865
rect 76146 275141 76346 275151
rect 76146 274961 76156 275141
rect 76336 274961 76346 275141
rect 76146 274951 76346 274961
rect 76601 271042 77001 284196
rect 77400 283324 77800 296486
rect 77400 283144 77414 283324
rect 77786 283144 77800 283324
rect 77118 273990 77318 274000
rect 77118 273810 77128 273990
rect 77308 273810 77318 273990
rect 77118 273800 77318 273810
rect 76601 270862 76615 271042
rect 76987 270862 77001 271042
rect 76157 264562 76357 264572
rect 76157 264382 76167 264562
rect 76347 264382 76357 264562
rect 76157 264372 76357 264382
rect 55321 263511 75955 263611
rect 55321 57706 55421 263511
rect 76169 261803 76369 261813
rect 76169 261623 76179 261803
rect 76359 261623 76369 261803
rect 76169 261613 76369 261623
rect 76601 257698 77001 270862
rect 77400 269977 77800 283144
rect 77400 269797 77414 269977
rect 77786 269797 77800 269977
rect 77120 260645 77320 260655
rect 77120 260465 77130 260645
rect 77310 260465 77320 260645
rect 77120 260455 77320 260465
rect 76601 257518 76615 257698
rect 76987 257518 77001 257698
rect 76154 251213 76354 251223
rect 76154 251033 76164 251213
rect 76344 251033 76354 251213
rect 76154 251023 76354 251033
rect 55759 250170 75947 250270
rect 55759 58068 55859 250170
rect 76152 248454 76352 248464
rect 76152 248274 76162 248454
rect 76342 248274 76352 248454
rect 76152 248264 76352 248274
rect 76601 244362 77001 257518
rect 77400 256634 77800 269797
rect 77400 256454 77414 256634
rect 77786 256454 77800 256634
rect 77098 247298 77298 247308
rect 77098 247118 77108 247298
rect 77288 247118 77298 247298
rect 77098 247108 77298 247118
rect 76601 244352 77002 244362
rect 76601 244172 76616 244352
rect 76988 244172 77002 244352
rect 76601 244162 77002 244172
rect 76201 237840 76401 237850
rect 76201 237660 76211 237840
rect 76391 237660 76401 237840
rect 76201 237650 76401 237660
rect 56349 236795 76055 236895
rect 56349 58593 56449 236795
rect 76199 235072 76399 235082
rect 76199 234892 76209 235072
rect 76389 234892 76399 235072
rect 76199 234882 76399 234892
rect 76601 230979 77001 244162
rect 77400 243289 77800 256454
rect 77400 243109 77414 243289
rect 77786 243109 77800 243289
rect 77076 233916 77276 233926
rect 77076 233736 77086 233916
rect 77266 233736 77276 233916
rect 77076 233726 77276 233736
rect 76601 230969 77003 230979
rect 76601 230789 76617 230969
rect 76989 230789 77003 230969
rect 76601 230779 77003 230789
rect 76601 216543 77001 230779
rect 76601 216167 76613 216543
rect 76989 216167 77001 216543
rect 76601 213299 77001 216167
rect 77400 229910 77800 243109
rect 77400 229730 77414 229910
rect 77786 229730 77800 229910
rect 77400 215798 77800 229730
rect 78409 322048 78809 335203
rect 79433 333954 79833 347097
rect 79433 333944 79835 333954
rect 79433 333764 79449 333944
rect 79821 333764 79835 333944
rect 79433 333754 79835 333764
rect 79011 326420 79211 326430
rect 79011 326240 79021 326420
rect 79201 326240 79211 326420
rect 79011 326230 79211 326240
rect 78409 321868 78423 322048
rect 78795 321868 78809 322048
rect 78409 308713 78809 321868
rect 79433 320606 79833 333754
rect 79433 320596 79838 320606
rect 79433 320416 79452 320596
rect 79824 320416 79838 320596
rect 79433 320406 79838 320416
rect 78970 313082 79170 313092
rect 78970 312902 78980 313082
rect 79160 312902 79170 313082
rect 78970 312892 79170 312902
rect 78409 308703 78810 308713
rect 78409 308523 78424 308703
rect 78796 308523 78810 308703
rect 78409 308513 78810 308523
rect 78409 295368 78809 308513
rect 79433 307261 79833 320406
rect 79431 307251 79833 307261
rect 79431 307071 79445 307251
rect 79817 307071 79833 307251
rect 79431 307061 79833 307071
rect 78983 299731 79183 299741
rect 78983 299551 78993 299731
rect 79173 299551 79183 299731
rect 78983 299541 79183 299551
rect 78409 295358 78811 295368
rect 78409 295178 78425 295358
rect 78797 295178 78811 295358
rect 78409 295168 78811 295178
rect 78409 282013 78809 295168
rect 79433 293916 79833 307061
rect 79433 293906 79837 293916
rect 79433 293726 79451 293906
rect 79823 293726 79837 293906
rect 79433 293716 79837 293726
rect 78981 286388 79181 286398
rect 78981 286208 78991 286388
rect 79171 286208 79181 286388
rect 78981 286198 79181 286208
rect 78409 281833 78423 282013
rect 78795 281833 78809 282013
rect 78409 268683 78809 281833
rect 79433 280568 79833 293716
rect 79433 280388 79447 280568
rect 79819 280388 79833 280568
rect 78988 273049 79188 273059
rect 78988 272869 78998 273049
rect 79178 272869 79188 273049
rect 78988 272859 79188 272869
rect 78409 268673 78810 268683
rect 78409 268493 78424 268673
rect 78796 268493 78810 268673
rect 78409 268483 78810 268493
rect 78409 255323 78809 268483
rect 79433 267225 79833 280388
rect 79433 267215 79836 267225
rect 79433 267035 79450 267215
rect 79822 267035 79836 267215
rect 79433 267025 79836 267035
rect 78975 259698 79175 259708
rect 78975 259518 78985 259698
rect 79165 259518 79175 259698
rect 78975 259508 79175 259518
rect 78409 255143 78423 255323
rect 78795 255143 78809 255323
rect 78409 241983 78809 255143
rect 79433 253886 79833 267025
rect 121307 254790 121507 254800
rect 121307 254610 121317 254790
rect 121497 254610 121507 254790
rect 121307 254600 121507 254610
rect 79433 253876 79836 253886
rect 79433 253696 79450 253876
rect 79822 253696 79836 253876
rect 79433 253686 79836 253696
rect 78989 246352 79189 246362
rect 78989 246172 78999 246352
rect 79179 246172 79189 246352
rect 78989 246162 79189 246172
rect 78409 241973 78811 241983
rect 78409 241793 78425 241973
rect 78797 241793 78811 241973
rect 78409 241783 78811 241793
rect 78409 228609 78809 241783
rect 79433 240538 79833 253686
rect 79433 240528 79837 240538
rect 79433 240348 79451 240528
rect 79823 240348 79837 240528
rect 79433 240338 79837 240348
rect 78984 232970 79184 232980
rect 78984 232790 78994 232970
rect 79174 232790 79184 232970
rect 78984 232780 79184 232790
rect 78407 228599 78809 228609
rect 78407 228419 78421 228599
rect 78793 228419 78809 228599
rect 78407 228409 78809 228419
rect 77399 215786 77800 215798
rect 77399 215410 77411 215786
rect 77787 215410 77800 215786
rect 77399 215398 77800 215410
rect 77400 213297 77800 215398
rect 78409 214918 78809 228409
rect 79433 227157 79833 240338
rect 79431 227147 79833 227157
rect 79431 226967 79445 227147
rect 79817 226967 79833 227147
rect 79431 226957 79833 226967
rect 78409 214906 78810 214918
rect 78409 214530 78422 214906
rect 78798 214530 78810 214906
rect 78409 214518 78810 214530
rect 78409 213338 78809 214518
rect 79433 214128 79833 226957
rect 96730 225136 96930 225168
rect 96730 225000 96762 225136
rect 96898 225000 96930 225136
rect 96730 224968 96930 225000
rect 221701 216555 221901 216557
rect 310997 216555 311197 216557
rect 362298 216555 362498 216556
rect 452556 216555 452756 216563
rect 81977 216549 490752 216555
rect 81977 216543 452566 216549
rect 81977 216542 221711 216543
rect 81977 216166 82023 216542
rect 82399 216541 221711 216542
rect 82399 216540 208407 216541
rect 82399 216539 119112 216540
rect 82399 216167 93801 216539
rect 93981 216538 119112 216539
rect 93981 216167 106151 216538
rect 82399 216166 106151 216167
rect 106331 216168 119112 216538
rect 119292 216539 196063 216540
rect 119292 216538 182755 216539
rect 119292 216168 131456 216538
rect 106331 216166 131456 216168
rect 131636 216537 157106 216538
rect 131636 216166 144763 216537
rect 81977 216165 144763 216166
rect 144943 216166 157106 216537
rect 157286 216166 170408 216538
rect 170588 216167 182755 216538
rect 182935 216168 196063 216539
rect 196243 216169 208407 216540
rect 208587 216171 221711 216541
rect 221891 216541 311007 216543
rect 221891 216171 234062 216541
rect 208587 216169 234062 216171
rect 234242 216540 259712 216541
rect 234242 216169 247363 216540
rect 196243 216168 247363 216169
rect 247543 216169 259712 216540
rect 259892 216539 298660 216541
rect 259892 216534 285357 216539
rect 259892 216169 273011 216534
rect 247543 216168 273011 216169
rect 182935 216167 273011 216168
rect 170588 216166 273011 216167
rect 144943 216165 273011 216166
rect 81977 216162 273011 216165
rect 273191 216167 285357 216534
rect 285537 216169 298660 216539
rect 298840 216171 311007 216541
rect 311187 216542 452566 216543
rect 311187 216540 362308 216542
rect 311187 216534 336657 216540
rect 311187 216171 324312 216534
rect 298840 216169 324312 216171
rect 285537 216167 324312 216169
rect 273191 216162 324312 216167
rect 324492 216168 336657 216534
rect 336837 216538 362308 216540
rect 336837 216168 349963 216538
rect 324492 216166 349963 216168
rect 350143 216170 362308 216538
rect 362488 216540 452566 216542
rect 362488 216539 439256 216540
rect 362488 216538 426912 216539
rect 362488 216537 413612 216538
rect 362488 216534 401262 216537
rect 362488 216170 375606 216534
rect 350143 216166 375606 216170
rect 324492 216162 375606 216166
rect 375786 216162 387955 216534
rect 388135 216165 401262 216534
rect 401442 216166 413612 216537
rect 413792 216167 426912 216538
rect 427092 216168 439256 216539
rect 439436 216177 452566 216540
rect 452746 216541 490752 216549
rect 452746 216539 478211 216541
rect 452746 216177 464906 216539
rect 439436 216168 464906 216177
rect 427092 216167 464906 216168
rect 465086 216169 478211 216539
rect 478391 216535 490752 216541
rect 478391 216169 490553 216535
rect 465086 216167 490553 216169
rect 413792 216166 490553 216167
rect 401442 216165 490553 216166
rect 388135 216163 490553 216165
rect 490733 216163 490752 216535
rect 388135 216162 490752 216163
rect 81977 216155 490752 216162
rect 82011 216154 82411 216155
rect 93791 216153 93991 216155
rect 106141 216152 106341 216155
rect 119102 216154 119302 216155
rect 131446 216152 131646 216155
rect 144753 216151 144953 216155
rect 157096 216152 157296 216155
rect 170398 216152 170598 216155
rect 182745 216153 182945 216155
rect 196053 216154 196253 216155
rect 247353 216154 247553 216155
rect 273001 216148 273201 216155
rect 285347 216153 285547 216155
rect 324302 216148 324502 216155
rect 336647 216154 336847 216155
rect 349953 216152 350153 216155
rect 375596 216148 375796 216155
rect 387945 216148 388145 216155
rect 401252 216151 401452 216155
rect 413602 216152 413802 216155
rect 426902 216153 427102 216155
rect 439246 216154 439446 216155
rect 464896 216153 465096 216155
rect 490543 216149 490743 216155
rect 197110 215799 197310 215800
rect 209458 215799 209658 215800
rect 222764 215799 222964 215800
rect 235107 215799 235307 215800
rect 260760 215799 260960 215800
rect 299709 215799 299909 215800
rect 312056 215799 312256 215800
rect 389004 215799 389204 215801
rect 427961 215799 428161 215802
rect 453612 215799 453812 215802
rect 465958 215799 466158 215800
rect 82007 215788 491813 215799
rect 82007 215787 427971 215788
rect 82007 215411 82026 215787
rect 82402 215786 389014 215787
rect 82402 215785 197120 215786
rect 82402 215413 94858 215785
rect 95038 215413 107208 215785
rect 107388 215413 120173 215785
rect 120353 215782 145824 215785
rect 120353 215413 132517 215782
rect 82402 215411 132517 215413
rect 82007 215410 132517 215411
rect 132697 215413 145824 215782
rect 146004 215784 183817 215785
rect 146004 215778 171474 215784
rect 146004 215413 158164 215778
rect 132697 215410 158164 215413
rect 82007 215406 158164 215410
rect 158344 215412 171474 215778
rect 171654 215413 183817 215784
rect 183997 215414 197120 215785
rect 197300 215414 209468 215786
rect 209648 215414 222774 215786
rect 222954 215414 235117 215786
rect 235297 215785 260770 215786
rect 235297 215414 248419 215785
rect 183997 215413 248419 215414
rect 248599 215414 260770 215785
rect 260950 215784 299719 215786
rect 260950 215414 274071 215784
rect 248599 215413 274071 215414
rect 171654 215412 274071 215413
rect 274251 215412 286415 215784
rect 286595 215414 299719 215784
rect 299899 215414 312066 215786
rect 312246 215784 389014 215786
rect 312246 215414 325371 215784
rect 286595 215412 325371 215414
rect 325551 215781 351018 215784
rect 325551 215412 337716 215781
rect 158344 215409 337716 215412
rect 337896 215412 351018 215781
rect 351198 215412 363367 215784
rect 363547 215781 389014 215784
rect 363547 215412 376672 215781
rect 337896 215409 376672 215412
rect 376852 215415 389014 215781
rect 389194 215783 427971 215787
rect 389194 215415 402321 215783
rect 376852 215411 402321 215415
rect 402501 215781 427971 215783
rect 402501 215411 414668 215781
rect 376852 215409 414668 215411
rect 414848 215416 427971 215781
rect 428151 215782 453622 215788
rect 428151 215416 440316 215782
rect 414848 215410 440316 215416
rect 440496 215416 453622 215782
rect 453802 215786 491813 215788
rect 453802 215416 465968 215786
rect 440496 215414 465968 215416
rect 466148 215784 491813 215786
rect 466148 215414 479269 215784
rect 440496 215412 479269 215414
rect 479449 215412 491616 215784
rect 491796 215412 491813 215784
rect 440496 215410 491813 215412
rect 414848 215409 491813 215410
rect 158344 215406 491813 215409
rect 82007 215399 491813 215406
rect 132507 215396 132707 215399
rect 158154 215392 158354 215399
rect 171464 215398 171664 215399
rect 274061 215398 274261 215399
rect 286405 215398 286605 215399
rect 325361 215398 325561 215399
rect 337706 215395 337906 215399
rect 351008 215398 351208 215399
rect 363357 215398 363557 215399
rect 376662 215395 376862 215399
rect 402311 215397 402511 215399
rect 414658 215395 414858 215399
rect 440306 215396 440506 215399
rect 479259 215398 479459 215399
rect 491606 215398 491806 215399
rect 257695 215290 257895 215300
rect 232046 215275 232246 215285
rect 117109 215263 117309 215273
rect 91790 215250 91990 215260
rect 91790 215070 91800 215250
rect 91980 215070 91990 215250
rect 91790 215060 91990 215070
rect 104135 215241 104335 215251
rect 104135 215061 104145 215241
rect 104325 215061 104335 215241
rect 117109 215083 117119 215263
rect 117299 215083 117309 215263
rect 194044 215263 194244 215273
rect 155099 215247 155299 215257
rect 142759 215217 142959 215227
rect 117109 215073 117309 215083
rect 129444 215201 129644 215211
rect 104135 215051 104335 215061
rect 129444 215021 129454 215201
rect 129634 215021 129644 215201
rect 142759 215037 142769 215217
rect 142949 215037 142959 215217
rect 155099 215067 155109 215247
rect 155289 215067 155299 215247
rect 180755 215235 180955 215245
rect 155099 215057 155299 215067
rect 168401 215204 168601 215214
rect 142759 215027 142959 215037
rect 129444 215011 129644 215021
rect 168401 215024 168411 215204
rect 168591 215024 168601 215204
rect 180755 215055 180765 215235
rect 180945 215055 180955 215235
rect 194044 215083 194054 215263
rect 194234 215083 194244 215263
rect 194044 215073 194244 215083
rect 206402 215241 206602 215251
rect 180755 215045 180955 215055
rect 206402 215061 206412 215241
rect 206592 215061 206602 215241
rect 206402 215051 206602 215061
rect 219699 215240 219899 215250
rect 219699 215060 219709 215240
rect 219889 215060 219899 215240
rect 232046 215095 232056 215275
rect 232236 215095 232246 215275
rect 232046 215085 232246 215095
rect 245350 215259 245550 215269
rect 245350 215079 245360 215259
rect 245540 215079 245550 215259
rect 257695 215110 257705 215290
rect 257885 215110 257895 215290
rect 257695 215100 257895 215110
rect 271004 215271 271204 215281
rect 271004 215091 271014 215271
rect 271194 215091 271204 215271
rect 271004 215081 271204 215091
rect 283347 215253 283547 215263
rect 245350 215069 245550 215079
rect 283347 215073 283357 215253
rect 283537 215073 283547 215253
rect 283347 215063 283547 215073
rect 296650 215249 296850 215259
rect 296650 215069 296660 215249
rect 296840 215069 296850 215249
rect 219699 215050 219899 215060
rect 296650 215059 296850 215069
rect 308994 215256 309194 215266
rect 308994 215076 309004 215256
rect 309184 215076 309194 215256
rect 334645 215263 334845 215273
rect 308994 215066 309194 215076
rect 322301 215233 322501 215243
rect 322301 215053 322311 215233
rect 322491 215053 322501 215233
rect 334645 215083 334655 215263
rect 334835 215083 334845 215263
rect 385945 215264 386145 215274
rect 360295 215245 360495 215255
rect 334645 215073 334845 215083
rect 347951 215233 348151 215243
rect 322301 215043 322501 215053
rect 347951 215053 347961 215233
rect 348141 215053 348151 215233
rect 360295 215065 360305 215245
rect 360485 215065 360495 215245
rect 360295 215055 360495 215065
rect 373600 215237 373800 215247
rect 373600 215057 373610 215237
rect 373790 215057 373800 215237
rect 385945 215084 385955 215264
rect 386135 215084 386145 215264
rect 385945 215074 386145 215084
rect 399250 215263 399450 215273
rect 399250 215083 399260 215263
rect 399440 215083 399450 215263
rect 437247 215250 437447 215260
rect 399250 215073 399450 215083
rect 411599 215229 411799 215239
rect 347951 215043 348151 215053
rect 373600 215047 373800 215057
rect 411599 215049 411609 215229
rect 411789 215049 411799 215229
rect 411599 215039 411799 215049
rect 424899 215232 425099 215242
rect 424899 215052 424909 215232
rect 425089 215052 425099 215232
rect 437247 215070 437257 215250
rect 437437 215070 437447 215250
rect 437247 215060 437447 215070
rect 450543 215250 450743 215260
rect 450543 215070 450553 215250
rect 450733 215070 450743 215250
rect 450543 215060 450743 215070
rect 462894 215237 463094 215247
rect 424899 215042 425099 215052
rect 462894 215057 462904 215237
rect 463084 215057 463094 215237
rect 488547 215243 488747 215253
rect 462894 215047 463094 215057
rect 476206 215225 476406 215235
rect 476206 215045 476216 215225
rect 476396 215045 476406 215225
rect 488547 215063 488557 215243
rect 488737 215063 488747 215243
rect 488547 215053 488747 215063
rect 476206 215035 476406 215045
rect 168401 215014 168601 215024
rect 96165 214917 96365 214918
rect 108508 214917 108708 214921
rect 159470 214917 159670 214920
rect 172774 214917 172974 214918
rect 185121 214917 185321 214918
rect 224078 214917 224278 214920
rect 236418 214917 236618 214918
rect 262070 214917 262270 214919
rect 301030 214917 301230 214920
rect 313368 214917 313568 214918
rect 339018 214917 339218 214918
rect 364669 214917 364869 214918
rect 377974 214917 378174 214918
rect 441618 214917 441818 214918
rect 454924 214917 455124 214921
rect 82007 214907 493126 214917
rect 82007 214905 108518 214907
rect 82007 214529 82044 214905
rect 82420 214904 108518 214905
rect 82420 214532 96175 214904
rect 96355 214535 108518 214904
rect 108698 214906 454934 214907
rect 108698 214903 159480 214906
rect 108698 214901 133828 214903
rect 108698 214535 121484 214901
rect 96355 214532 121484 214535
rect 82420 214529 121484 214532
rect 121664 214531 133828 214901
rect 134008 214531 147132 214903
rect 147312 214534 159480 214903
rect 159660 214904 224088 214906
rect 159660 214534 172784 214904
rect 147312 214532 172784 214534
rect 172964 214532 185131 214904
rect 185311 214903 224088 214904
rect 185311 214902 210781 214903
rect 185311 214532 198432 214902
rect 147312 214531 198432 214532
rect 121664 214530 198432 214531
rect 198612 214531 210781 214902
rect 210961 214534 224088 214903
rect 224268 214905 301040 214906
rect 224268 214904 262080 214905
rect 224268 214534 236428 214904
rect 210961 214532 236428 214534
rect 236608 214901 262080 214904
rect 236608 214532 249732 214901
rect 210961 214531 249732 214532
rect 198612 214530 249732 214531
rect 121664 214529 249732 214530
rect 249912 214533 262080 214901
rect 262260 214903 301040 214905
rect 262260 214533 275383 214903
rect 249912 214531 275383 214533
rect 275563 214531 287731 214903
rect 287911 214534 301040 214903
rect 301220 214904 454934 214906
rect 301220 214534 313378 214904
rect 287911 214532 313378 214534
rect 313558 214903 339028 214904
rect 313558 214532 326683 214903
rect 287911 214531 326683 214532
rect 326863 214532 339028 214903
rect 339208 214901 364679 214904
rect 339208 214532 352334 214901
rect 326863 214531 352334 214532
rect 249912 214529 352334 214531
rect 352514 214532 364679 214901
rect 364859 214532 377984 214904
rect 378164 214902 441628 214904
rect 378164 214532 390331 214902
rect 352514 214530 390331 214532
rect 390511 214901 441628 214902
rect 390511 214898 429286 214901
rect 390511 214894 415976 214898
rect 390511 214530 403624 214894
rect 352514 214529 403624 214530
rect 82007 214522 403624 214529
rect 403804 214526 415976 214894
rect 416156 214529 429286 214898
rect 429466 214532 441628 214901
rect 441808 214535 454934 214904
rect 455114 214902 493126 214907
rect 455114 214535 467278 214902
rect 441808 214532 467278 214535
rect 429466 214530 467278 214532
rect 467458 214901 492932 214902
rect 467458 214530 480579 214901
rect 429466 214529 480579 214530
rect 480759 214530 492932 214901
rect 493112 214530 493126 214902
rect 480759 214529 493126 214530
rect 416156 214526 493126 214529
rect 403804 214522 493126 214526
rect 82007 214517 493126 214522
rect 121474 214515 121674 214517
rect 198422 214516 198622 214517
rect 249722 214515 249922 214517
rect 352324 214515 352524 214517
rect 390321 214516 390521 214517
rect 403614 214508 403814 214517
rect 415966 214512 416166 214517
rect 429276 214515 429476 214517
rect 467268 214516 467468 214517
rect 480569 214515 480769 214517
rect 492922 214516 493122 214517
rect 186585 214130 186785 214137
rect 212226 214130 212426 214133
rect 263531 214130 263731 214134
rect 340473 214130 340673 214131
rect 366116 214130 366316 214132
rect 379434 214130 379634 214131
rect 417427 214130 417627 214134
rect 430742 214130 430942 214133
rect 468736 214130 468936 214133
rect 496671 214130 497071 549638
rect 79432 214116 79833 214128
rect 79432 213740 79444 214116
rect 79820 213740 79833 214116
rect 79432 213728 79833 213740
rect 82022 214123 497071 214130
rect 82022 214117 186595 214123
rect 82022 213741 82058 214117
rect 82434 214116 186595 214117
rect 82434 214115 122935 214116
rect 82434 213743 97623 214115
rect 97803 214111 122935 214115
rect 97803 213743 109981 214111
rect 82434 213741 109981 213743
rect 82022 213739 109981 213741
rect 110161 213744 122935 214111
rect 123115 214113 186595 214116
rect 123115 213744 135298 214113
rect 110161 213741 135298 213744
rect 135478 214111 186595 214113
rect 135478 214105 174235 214111
rect 135478 213741 148591 214105
rect 110161 213739 148591 213741
rect 82022 213733 148591 213739
rect 148771 213733 160931 214105
rect 161111 213739 174235 214105
rect 174415 213751 186595 214111
rect 186775 214120 497071 214123
rect 186775 214119 263541 214120
rect 186775 214105 212236 214119
rect 186775 213751 199887 214105
rect 174415 213739 199887 213751
rect 161111 213733 199887 213739
rect 200067 213747 212236 214105
rect 212416 214116 263541 214119
rect 212416 214115 251199 214116
rect 212416 214113 237896 214115
rect 212416 213747 225542 214113
rect 200067 213741 225542 213747
rect 225722 213743 237896 214113
rect 238076 213744 251199 214115
rect 251379 213748 263541 214116
rect 263721 214118 417437 214120
rect 263721 214117 366126 214118
rect 263721 214116 340483 214117
rect 263721 214113 314835 214116
rect 263721 214111 302496 214113
rect 263721 213748 276848 214111
rect 251379 213744 276848 213748
rect 238076 213743 276848 213744
rect 225722 213741 276848 213743
rect 200067 213739 276848 213741
rect 277028 214110 302496 214111
rect 277028 213739 289177 214110
rect 200067 213738 289177 213739
rect 289357 213741 302496 214110
rect 302676 213744 314835 214113
rect 315015 213744 328133 214116
rect 328313 213745 340483 214116
rect 340663 214113 366126 214117
rect 340663 213745 353792 214113
rect 328313 213744 353792 213745
rect 302676 213741 353792 213744
rect 353972 213746 366126 214113
rect 366306 214117 417437 214118
rect 366306 213746 379444 214117
rect 353972 213745 379444 213746
rect 379624 214114 417437 214117
rect 379624 213745 391778 214114
rect 353972 213742 391778 213745
rect 391958 214110 417437 214114
rect 391958 213742 405089 214110
rect 353972 213741 405089 213742
rect 289357 213738 405089 213741
rect 405269 213748 417437 214110
rect 417617 214119 497071 214120
rect 417617 213748 430752 214119
rect 405269 213747 430752 213748
rect 430932 214113 468746 214119
rect 430932 213747 443088 214113
rect 405269 213741 443088 213747
rect 443268 213741 456393 214113
rect 456573 213747 468746 214113
rect 468926 214114 497071 214119
rect 468926 214113 494383 214114
rect 468926 213747 482048 214113
rect 456573 213741 482048 213747
rect 482228 213742 494383 214113
rect 494563 213742 497071 214114
rect 482228 213741 497071 213742
rect 405269 213738 497071 213741
rect 200067 213733 497071 213738
rect 82022 213730 497071 213733
rect 82046 213729 82446 213730
rect 97613 213729 97813 213730
rect 79433 213416 79833 213728
rect 109971 213725 110171 213730
rect 135288 213727 135488 213730
rect 148581 213719 148781 213730
rect 160921 213719 161121 213730
rect 174225 213725 174425 213730
rect 199877 213719 200077 213730
rect 225532 213727 225732 213730
rect 237886 213729 238086 213730
rect 276838 213725 277038 213730
rect 289167 213724 289367 213730
rect 302486 213727 302686 213730
rect 353782 213727 353982 213730
rect 391768 213728 391968 213730
rect 405079 213724 405279 213730
rect 443078 213727 443278 213730
rect 456383 213727 456583 213730
rect 482038 213727 482238 213730
rect 494373 213728 494573 213730
rect 436200 213531 436600 213543
rect 90843 213445 91043 213455
rect 90843 213265 90853 213445
rect 91033 213265 91043 213445
rect 90843 213255 91043 213265
rect 103193 213443 103393 213453
rect 103193 213263 103203 213443
rect 103383 213263 103393 213443
rect 103193 213253 103393 213263
rect 116153 213444 116353 213454
rect 116153 213264 116163 213444
rect 116343 213264 116353 213444
rect 347002 213441 347202 213451
rect 154145 213428 154345 213438
rect 116153 213254 116353 213264
rect 128496 213403 128696 213413
rect 128496 213223 128506 213403
rect 128686 213223 128696 213403
rect 128496 213213 128696 213223
rect 141801 213363 142001 213373
rect 141801 213183 141811 213363
rect 141991 213183 142001 213363
rect 154145 213248 154155 213428
rect 154335 213248 154345 213428
rect 179800 213423 180000 213433
rect 205446 213429 205646 213439
rect 154145 213238 154345 213248
rect 167456 213389 167656 213399
rect 167456 213209 167466 213389
rect 167646 213209 167656 213389
rect 179800 213243 179810 213423
rect 179990 213243 180000 213423
rect 179800 213233 180000 213243
rect 193110 213415 193310 213425
rect 193110 213235 193120 213415
rect 193300 213235 193310 213415
rect 205446 213249 205456 213429
rect 205636 213249 205646 213429
rect 205446 213239 205646 213249
rect 218751 213430 218951 213440
rect 218751 213250 218761 213430
rect 218941 213250 218951 213430
rect 256749 213427 256949 213437
rect 218751 213240 218951 213250
rect 231101 213417 231301 213427
rect 193110 213225 193310 213235
rect 231101 213237 231111 213417
rect 231291 213237 231301 213417
rect 231101 213227 231301 213237
rect 244400 213407 244600 213417
rect 244400 213227 244410 213407
rect 244590 213227 244600 213407
rect 256749 213247 256759 213427
rect 256939 213247 256949 213427
rect 256749 213237 256949 213247
rect 270058 213408 270258 213418
rect 321351 213417 321551 213427
rect 244400 213217 244600 213227
rect 270058 213228 270068 213408
rect 270248 213228 270258 213408
rect 295705 213400 295905 213410
rect 270058 213218 270258 213228
rect 282402 213385 282602 213395
rect 167456 213199 167656 213209
rect 282402 213205 282412 213385
rect 282592 213205 282602 213385
rect 295705 213220 295715 213400
rect 295895 213220 295905 213400
rect 295705 213210 295905 213220
rect 308053 213358 308253 213368
rect 282402 213195 282602 213205
rect 141801 213173 142001 213183
rect 308053 213178 308063 213358
rect 308243 213178 308253 213358
rect 321351 213237 321361 213417
rect 321541 213237 321551 213417
rect 321351 213227 321551 213237
rect 333696 213374 333896 213384
rect 333696 213194 333706 213374
rect 333886 213194 333896 213374
rect 347002 213261 347012 213441
rect 347192 213261 347202 213441
rect 372654 213441 372854 213451
rect 347002 213251 347202 213261
rect 359351 213429 359551 213439
rect 359351 213249 359361 213429
rect 359541 213249 359551 213429
rect 372654 213261 372664 213441
rect 372844 213261 372854 213441
rect 372654 213251 372854 213261
rect 385001 213442 385201 213452
rect 385001 213262 385011 213442
rect 385191 213262 385201 213442
rect 385001 213252 385201 213262
rect 398298 213437 398498 213447
rect 398298 213257 398308 213437
rect 398488 213257 398498 213437
rect 359351 213239 359551 213249
rect 398298 213247 398498 213257
rect 410646 213437 410846 213447
rect 410646 213257 410656 213437
rect 410836 213257 410846 213437
rect 410646 213247 410846 213257
rect 423955 213440 424155 213450
rect 423955 213260 423965 213440
rect 424145 213260 424155 213440
rect 423955 213250 424155 213260
rect 333696 213184 333896 213194
rect 308053 213168 308253 213178
rect 436200 213155 436212 213531
rect 436588 213155 436600 213531
rect 449605 213433 449805 213443
rect 449605 213253 449615 213433
rect 449795 213253 449805 213433
rect 449605 213243 449805 213253
rect 461953 213431 462153 213441
rect 461953 213251 461963 213431
rect 462143 213251 462153 213431
rect 461953 213241 462153 213251
rect 475250 213426 475450 213436
rect 475250 213246 475260 213426
rect 475440 213246 475450 213426
rect 475250 213236 475450 213246
rect 487598 213400 487798 213410
rect 487598 213220 487608 213400
rect 487788 213220 487798 213400
rect 487598 213210 487798 213220
rect 436200 213143 436600 213155
rect 86929 212784 87129 212794
rect 86929 212604 86939 212784
rect 87119 212604 87129 212784
rect 115001 212793 115201 212803
rect 112234 212768 112434 212778
rect 86929 212594 87129 212604
rect 89691 212753 89891 212763
rect 89691 212573 89701 212753
rect 89881 212573 89891 212753
rect 102047 212758 102247 212768
rect 89691 212563 89891 212573
rect 99274 212733 99474 212743
rect 99274 212553 99284 212733
rect 99464 212553 99474 212733
rect 102047 212578 102057 212758
rect 102237 212578 102247 212758
rect 112234 212588 112244 212768
rect 112424 212588 112434 212768
rect 115001 212613 115011 212793
rect 115191 212613 115201 212793
rect 332544 212788 332744 212798
rect 115001 212603 115201 212613
rect 124573 212758 124773 212768
rect 140651 212765 140851 212775
rect 112234 212578 112434 212588
rect 124573 212578 124583 212758
rect 124763 212578 124773 212758
rect 102047 212568 102247 212578
rect 124573 212568 124773 212578
rect 127346 212749 127546 212759
rect 127346 212569 127356 212749
rect 127536 212569 127546 212749
rect 127346 212559 127546 212569
rect 137889 212745 138089 212755
rect 137889 212565 137899 212745
rect 138079 212565 138089 212745
rect 140651 212585 140661 212765
rect 140841 212585 140851 212765
rect 214834 212767 215034 212777
rect 201526 212747 201726 212757
rect 152989 212722 153189 212732
rect 140651 212575 140851 212585
rect 150231 212706 150431 212716
rect 137889 212555 138089 212565
rect 99274 212543 99474 212553
rect 150231 212526 150241 212706
rect 150421 212526 150431 212706
rect 152989 212542 152999 212722
rect 153179 212542 153189 212722
rect 152989 212532 153189 212542
rect 163531 212723 163731 212733
rect 163531 212543 163541 212723
rect 163721 212543 163731 212723
rect 175881 212730 176081 212740
rect 163531 212533 163731 212543
rect 166302 212711 166502 212721
rect 150231 212516 150431 212526
rect 166302 212531 166312 212711
rect 166492 212531 166502 212711
rect 175881 212550 175891 212730
rect 176071 212550 176081 212730
rect 189185 212737 189385 212747
rect 175881 212540 176081 212550
rect 178642 212711 178842 212721
rect 166302 212521 166502 212531
rect 178642 212531 178652 212711
rect 178832 212531 178842 212711
rect 189185 212557 189195 212737
rect 189375 212557 189385 212737
rect 189185 212547 189385 212557
rect 191952 212737 192152 212747
rect 191952 212557 191962 212737
rect 192142 212557 192152 212737
rect 201526 212567 201536 212747
rect 201716 212567 201726 212747
rect 201526 212557 201726 212567
rect 204292 212725 204492 212735
rect 191952 212547 192152 212557
rect 204292 212545 204302 212725
rect 204482 212545 204492 212725
rect 214834 212587 214844 212767
rect 215024 212587 215034 212767
rect 214834 212577 215034 212587
rect 217598 212763 217798 212773
rect 217598 212583 217608 212763
rect 217788 212583 217798 212763
rect 217598 212573 217798 212583
rect 227185 212756 227385 212766
rect 227185 212576 227195 212756
rect 227375 212576 227385 212756
rect 240486 212755 240686 212765
rect 227185 212566 227385 212576
rect 229944 212734 230144 212744
rect 204292 212535 204492 212545
rect 229944 212554 229954 212734
rect 230134 212554 230144 212734
rect 240486 212575 240496 212755
rect 240676 212575 240686 212755
rect 240486 212565 240686 212575
rect 243247 212764 243447 212774
rect 243247 212584 243257 212764
rect 243437 212584 243447 212764
rect 243247 212574 243447 212584
rect 252832 212745 253032 212755
rect 252832 212565 252842 212745
rect 253022 212565 253032 212745
rect 252832 212555 253032 212565
rect 255592 212745 255792 212755
rect 329781 212753 329981 212763
rect 255592 212565 255602 212745
rect 255782 212565 255792 212745
rect 281245 212736 281445 212746
rect 278477 212726 278677 212736
rect 268900 212695 269100 212705
rect 255592 212555 255792 212565
rect 266133 212661 266333 212671
rect 229944 212544 230144 212554
rect 178642 212521 178842 212531
rect 266133 212481 266143 212661
rect 266323 212481 266333 212661
rect 268900 212515 268910 212695
rect 269090 212515 269100 212695
rect 278477 212546 278487 212726
rect 278667 212546 278677 212726
rect 281245 212556 281255 212736
rect 281435 212556 281445 212736
rect 317440 212726 317640 212736
rect 304137 212711 304337 212721
rect 294548 212691 294748 212701
rect 281245 212546 281445 212556
rect 291785 212670 291985 212680
rect 278477 212536 278677 212546
rect 268900 212505 269100 212515
rect 266133 212471 266333 212481
rect 291785 212490 291795 212670
rect 291975 212490 291985 212670
rect 294548 212511 294558 212691
rect 294738 212511 294748 212691
rect 304137 212531 304147 212711
rect 304327 212531 304337 212711
rect 304137 212521 304337 212531
rect 306901 212706 307101 212716
rect 306901 212526 306911 212706
rect 307091 212526 307101 212706
rect 317440 212546 317450 212726
rect 317630 212546 317640 212726
rect 317440 212536 317640 212546
rect 320198 212726 320398 212736
rect 320198 212546 320208 212726
rect 320388 212546 320398 212726
rect 329781 212573 329791 212753
rect 329971 212573 329981 212753
rect 332544 212608 332554 212788
rect 332734 212608 332744 212788
rect 383846 212772 384046 212782
rect 381081 212753 381281 212763
rect 358194 212739 358394 212749
rect 332544 212598 332744 212608
rect 343087 212724 343287 212734
rect 329781 212563 329981 212573
rect 320198 212536 320398 212546
rect 343087 212544 343097 212724
rect 343277 212544 343287 212724
rect 343087 212534 343287 212544
rect 345849 212729 346049 212739
rect 345849 212549 345859 212729
rect 346039 212549 346049 212729
rect 345849 212539 346049 212549
rect 355428 212720 355628 212730
rect 355428 212540 355438 212720
rect 355618 212540 355628 212720
rect 358194 212559 358204 212739
rect 358384 212559 358394 212739
rect 371499 212730 371699 212740
rect 358194 212549 358394 212559
rect 368737 212706 368937 212716
rect 355428 212530 355628 212540
rect 306901 212516 307101 212526
rect 368737 212526 368747 212706
rect 368927 212526 368937 212706
rect 371499 212550 371509 212730
rect 371689 212550 371699 212730
rect 381081 212573 381091 212753
rect 381271 212573 381281 212753
rect 383846 212592 383856 212772
rect 384036 212592 384046 212772
rect 397149 212767 397349 212777
rect 422800 212776 423000 212786
rect 383846 212582 384046 212592
rect 394388 212717 394588 212727
rect 381081 212563 381281 212573
rect 371499 212540 371699 212550
rect 394388 212537 394398 212717
rect 394578 212537 394588 212717
rect 397149 212587 397159 212767
rect 397339 212587 397349 212767
rect 409496 212753 409696 212763
rect 397149 212577 397349 212587
rect 406727 212733 406927 212743
rect 406727 212553 406737 212733
rect 406917 212553 406927 212733
rect 409496 212573 409506 212753
rect 409686 212573 409696 212753
rect 409496 212563 409696 212573
rect 420037 212758 420237 212768
rect 420037 212578 420047 212758
rect 420227 212578 420237 212758
rect 422800 212596 422810 212776
rect 422990 212596 423000 212776
rect 422800 212586 423000 212596
rect 432386 212773 432586 212783
rect 432386 212593 432396 212773
rect 432576 212593 432586 212773
rect 432386 212583 432586 212593
rect 435145 212745 435345 212755
rect 420037 212568 420237 212578
rect 435145 212565 435155 212745
rect 435335 212565 435345 212745
rect 448449 212744 448649 212754
rect 435145 212555 435345 212565
rect 445681 212690 445881 212700
rect 406727 212543 406927 212553
rect 394388 212527 394588 212537
rect 368737 212516 368937 212526
rect 294548 212501 294748 212511
rect 445681 212510 445691 212690
rect 445871 212510 445881 212690
rect 448449 212564 448459 212744
rect 448639 212564 448649 212744
rect 460793 212737 460993 212747
rect 448449 212554 448649 212564
rect 458031 212705 458231 212715
rect 458031 212525 458041 212705
rect 458221 212525 458231 212705
rect 460793 212557 460803 212737
rect 460983 212557 460993 212737
rect 486447 212741 486647 212751
rect 474100 212713 474300 212723
rect 460793 212547 460993 212557
rect 471328 212659 471528 212669
rect 458031 212515 458231 212525
rect 445681 212500 445881 212510
rect 291785 212480 291985 212490
rect 471328 212479 471338 212659
rect 471518 212479 471528 212659
rect 474100 212533 474110 212713
rect 474290 212533 474300 212713
rect 474100 212523 474300 212533
rect 483684 212671 483884 212681
rect 483684 212491 483694 212671
rect 483874 212491 483884 212671
rect 486447 212561 486457 212741
rect 486637 212561 486647 212741
rect 486447 212551 486647 212561
rect 483684 212481 483884 212491
rect 471328 212469 471528 212479
rect 101200 212328 101300 212350
rect 101200 212272 101222 212328
rect 101278 212272 101300 212328
rect 88853 191898 88953 212270
rect 100236 192094 100336 212260
rect 101200 212250 101300 212272
rect 126513 212315 126613 212337
rect 126513 212259 126535 212315
rect 126591 212259 126613 212315
rect 152164 212314 152264 212336
rect 100236 192038 100258 192094
rect 100314 192038 100336 192094
rect 100236 192016 100336 192038
rect 76286 191798 88953 191898
rect 76286 80900 76386 191798
rect 114150 190150 114250 212250
rect 125540 191953 125640 212254
rect 126513 212237 126613 212259
rect 125540 191931 125641 191953
rect 125540 191875 125563 191931
rect 125619 191875 125641 191931
rect 125540 191853 125641 191875
rect 77951 190050 114250 190150
rect 77951 82694 78051 190050
rect 139807 187581 139907 212305
rect 152164 212258 152186 212314
rect 152242 212258 152264 212314
rect 177803 212310 177903 212332
rect 152164 212236 152264 212258
rect 151197 189955 151297 212232
rect 151197 189899 151219 189955
rect 151275 189899 151297 189955
rect 151197 189877 151297 189899
rect 79033 187481 139907 187581
rect 79033 84107 79133 187481
rect 165463 184606 165563 212298
rect 176840 190325 176940 212275
rect 177803 212254 177825 212310
rect 177881 212254 177903 212310
rect 203459 212316 203559 212338
rect 177803 212232 177903 212254
rect 176840 190269 176862 190325
rect 176918 190269 176940 190325
rect 176840 190240 176940 190269
rect 80012 184506 165563 184606
rect 80012 85005 80112 184506
rect 191099 180979 191199 212262
rect 202478 188135 202578 212275
rect 203459 212260 203481 212316
rect 203537 212260 203559 212316
rect 229098 212316 229198 212338
rect 203459 212238 203559 212260
rect 202478 188113 202579 188135
rect 202478 188057 202501 188113
rect 202557 188057 202579 188113
rect 202478 188035 202579 188057
rect 202478 188027 202578 188035
rect 80949 180879 191199 180979
rect 80949 85436 81049 180879
rect 216743 178077 216843 212270
rect 228146 187406 228246 212268
rect 229098 212260 229120 212316
rect 229176 212260 229198 212316
rect 254765 212313 254865 212335
rect 229098 212238 229198 212260
rect 228146 187350 228168 187406
rect 228224 187350 228246 187406
rect 228146 187303 228246 187350
rect 81740 177977 216843 178077
rect 81740 85861 81840 177977
rect 242423 173480 242523 212287
rect 254765 212257 254787 212313
rect 254843 212257 254865 212313
rect 280408 212316 280508 212338
rect 253784 188715 253884 212243
rect 254765 212235 254865 212257
rect 253784 188659 253806 188715
rect 253862 188659 253884 188715
rect 253784 187320 253884 188659
rect 82928 173380 242523 173480
rect 82928 86327 83028 173380
rect 268056 169952 268156 212294
rect 279438 186937 279538 212270
rect 280408 212260 280430 212316
rect 280486 212260 280508 212316
rect 306061 212311 306161 212333
rect 280408 212238 280508 212260
rect 279438 186881 279460 186937
rect 279516 186881 279538 186937
rect 279438 186829 279538 186881
rect 83688 169852 268156 169952
rect 83688 86685 83788 169852
rect 293694 166499 293794 212264
rect 306061 212255 306083 212311
rect 306139 212255 306161 212311
rect 331707 212311 331807 212333
rect 305089 186372 305189 212252
rect 306061 212233 306161 212255
rect 305089 186316 305111 186372
rect 305167 186316 305189 186372
rect 305089 186287 305189 186316
rect 84369 166399 293794 166499
rect 84369 87093 84469 166399
rect 319341 162698 319441 212264
rect 330739 187409 330839 212281
rect 331707 212255 331729 212311
rect 331785 212255 331807 212311
rect 357354 212320 357454 212342
rect 331707 212233 331807 212255
rect 330739 187353 330761 187409
rect 330817 187353 330839 187409
rect 330739 187320 330839 187353
rect 85885 162598 319441 162698
rect 85885 87853 85985 162598
rect 344989 159544 345089 212279
rect 357354 212264 357376 212320
rect 357432 212264 357454 212320
rect 382989 212316 383089 212338
rect 356393 189652 356493 212254
rect 357354 212242 357454 212264
rect 356393 189596 356415 189652
rect 356471 189596 356493 189652
rect 356393 189557 356493 189596
rect 87620 159444 345089 159544
rect 87620 88461 87720 159444
rect 370673 157374 370773 212278
rect 382989 212260 383011 212316
rect 383067 212260 383089 212316
rect 408655 212316 408755 212338
rect 382031 191030 382131 212253
rect 382989 212238 383089 212260
rect 382031 190974 382053 191030
rect 382109 190974 382131 191030
rect 382031 190952 382131 190974
rect 88982 157274 370773 157374
rect 88982 89104 89082 157274
rect 396312 155153 396412 212254
rect 407703 192377 407803 212266
rect 408655 212260 408677 212316
rect 408733 212260 408755 212316
rect 434292 212311 434392 212333
rect 408655 212238 408755 212260
rect 407703 192321 407725 192377
rect 407781 192321 407803 192377
rect 407703 192297 407803 192321
rect 89997 155053 396412 155153
rect 89997 89570 90097 155053
rect 421951 151716 422051 212274
rect 433348 194511 433448 212260
rect 434292 212255 434314 212311
rect 434370 212255 434392 212311
rect 459957 212312 460057 212334
rect 434292 212233 434392 212255
rect 433348 194455 433370 194511
rect 433426 194455 433448 194511
rect 433348 194404 433448 194455
rect 90459 151616 422051 151716
rect 90459 89856 90559 151616
rect 447623 150035 447723 212278
rect 459957 212256 459979 212312
rect 460035 212256 460057 212312
rect 485598 212314 485698 212336
rect 458989 195926 459089 212237
rect 459957 212234 460057 212256
rect 458989 195870 459011 195926
rect 459067 195870 459089 195926
rect 458989 195820 459089 195870
rect 92066 149935 447723 150035
rect 92066 90451 92166 149935
rect 473285 145142 473385 212264
rect 485598 212258 485620 212314
rect 485676 212258 485698 212314
rect 484636 197100 484736 212252
rect 485598 212236 485698 212258
rect 484636 197044 484658 197100
rect 484714 197044 484736 197100
rect 484636 197017 484736 197044
rect 95014 145042 473385 145142
rect 95014 91512 95114 145042
rect 377541 103392 377741 103453
rect 377541 103336 377607 103392
rect 377663 103336 377741 103392
rect 373988 102680 374188 102742
rect 373988 102624 374062 102680
rect 374118 102624 374188 102680
rect 370445 101553 370645 101625
rect 370445 101497 370515 101553
rect 370571 101497 370645 101553
rect 366892 100538 367092 100599
rect 366892 100482 366968 100538
rect 367024 100482 367092 100538
rect 363354 99401 363554 99456
rect 363354 99345 363423 99401
rect 363479 99345 363554 99401
rect 359801 97974 360001 98044
rect 359801 97918 359877 97974
rect 359933 97918 360001 97974
rect 356258 95191 356458 95266
rect 356258 95135 356344 95191
rect 356400 95135 356458 95191
rect 352705 92852 352905 92937
rect 352705 92796 352774 92852
rect 352830 92796 352905 92852
rect 95014 91412 349373 91512
rect 92066 90402 345826 90451
rect 92066 90351 345827 90402
rect 90459 89756 342288 89856
rect 89997 89470 338741 89570
rect 88982 89004 335184 89104
rect 87620 88361 331638 88461
rect 85885 87753 328098 87853
rect 84369 86993 324552 87093
rect 83688 86684 321000 86685
rect 83688 86585 321002 86684
rect 82928 86230 317454 86327
rect 82928 86227 317455 86230
rect 81740 85761 313915 85861
rect 80949 85336 310369 85436
rect 80012 85004 306713 85005
rect 80012 84905 306812 85004
rect 79033 84007 303261 84107
rect 77951 82594 299726 82694
rect 76286 80700 296180 80900
rect 292436 78895 292636 78961
rect 292436 78843 292516 78895
rect 292568 78843 292636 78895
rect 288890 77835 289090 77894
rect 288890 77783 288955 77835
rect 289007 77783 289090 77835
rect 285350 76784 285550 76899
rect 285350 76732 285422 76784
rect 285474 76732 285550 76784
rect 281804 75137 282004 75240
rect 281804 75085 281872 75137
rect 281924 75085 282004 75137
rect 278247 74319 278447 74419
rect 278247 74267 278312 74319
rect 278364 74267 278447 74319
rect 274701 73242 274901 73381
rect 274701 73190 274773 73242
rect 274825 73190 274901 73242
rect 271161 71897 271361 72038
rect 271161 71845 271233 71897
rect 271285 71845 271361 71897
rect 267615 70521 267815 70588
rect 267615 70469 267693 70521
rect 267745 70469 267815 70521
rect 264065 69634 264265 69729
rect 264065 69582 264145 69634
rect 264197 69582 264265 69634
rect 260518 67282 260718 67416
rect 260518 67230 260593 67282
rect 260645 67230 260718 67282
rect 256978 66648 257178 66699
rect 256978 66596 257049 66648
rect 257101 66596 257178 66648
rect 253432 65352 253632 65406
rect 253432 65300 253511 65352
rect 253563 65300 253632 65352
rect 249875 64198 250075 64246
rect 249875 64146 249945 64198
rect 249997 64146 250075 64198
rect 246324 63355 246524 63441
rect 246324 63303 246384 63355
rect 246436 63303 246524 63355
rect 242789 62527 242989 62575
rect 242789 62475 242866 62527
rect 242918 62475 242989 62527
rect 239243 61793 239443 61871
rect 239243 61741 239313 61793
rect 239365 61741 239443 61793
rect 56349 58493 235901 58593
rect 55759 57968 232355 58068
rect 55321 57606 228815 57706
rect 54958 56648 225269 56748
rect 54700 56241 221712 56341
rect 54315 55957 218166 56057
rect 53978 55599 214626 55699
rect 53572 55075 211080 55175
rect 53197 54595 207530 54695
rect 52854 53882 203991 53982
rect 52556 53417 200443 53517
rect 52081 52370 196897 52470
rect 51598 51607 193340 51707
rect 50678 50868 189794 50968
rect 49956 49796 186254 49896
rect 48822 48594 182708 48694
rect 178966 46841 179166 46866
rect 178966 46789 179041 46841
rect 179093 46789 179166 46841
rect 175420 46565 175620 46590
rect 175420 46513 175484 46565
rect 175536 46513 175620 46565
rect 171880 46300 172080 46324
rect 171880 46248 171955 46300
rect 172007 46248 172080 46300
rect 168334 46061 168534 46094
rect 168334 46009 168401 46061
rect 168453 46009 168534 46061
rect 164777 45794 164977 45842
rect 164777 45742 164849 45794
rect 164901 45742 164977 45794
rect 161231 45504 161431 45566
rect 161231 45452 161304 45504
rect 161356 45452 161431 45504
rect 157691 45328 157891 45376
rect 157691 45276 157763 45328
rect 157815 45276 157891 45328
rect 154145 44976 154345 45073
rect 154145 44924 154216 44976
rect 154268 44924 154345 44976
rect 150595 44693 150795 44743
rect 150595 44641 150665 44693
rect 150717 44641 150795 44693
rect 147048 44470 147248 44527
rect 147048 44418 147097 44470
rect 147149 44418 147248 44470
rect 143508 44225 143708 44290
rect 143508 44173 143572 44225
rect 143624 44173 143708 44225
rect 139962 43855 140162 43905
rect 139962 43803 140048 43855
rect 140100 43803 140162 43855
rect 136405 43622 136605 43706
rect 136405 43570 136480 43622
rect 136532 43570 136605 43622
rect 132859 43380 133059 43419
rect 132859 43328 132931 43380
rect 132983 43328 133059 43380
rect 129319 43162 129519 43218
rect 129319 43110 129389 43162
rect 129441 43110 129519 43162
rect 125773 42860 125973 42920
rect 125773 42808 125856 42860
rect 125908 42808 125973 42860
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125773 363 125973 42808
rect 125816 -800 125928 363
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129319 326 129519 43110
rect 129362 -800 129474 326
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132859 221 133059 43328
rect 132908 -800 133020 221
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136405 11 136605 43570
rect 136454 -800 136566 11
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 139962 166 140162 43803
rect 140000 -800 140112 166
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143508 129 143708 44173
rect 143546 -800 143658 129
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147048 24 147248 44418
rect 147092 -800 147204 24
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150595 -6 150795 44641
rect 150638 -800 150750 -6
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154145 363 154345 44924
rect 154184 -800 154296 363
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157691 326 157891 45276
rect 157730 -800 157842 326
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161231 221 161431 45452
rect 161276 -800 161388 221
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164777 184 164977 45742
rect 164822 -800 164934 184
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168334 166 168534 46009
rect 168368 -800 168480 166
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171880 129 172080 46248
rect 171914 -800 172026 129
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175420 24 175620 46513
rect 175460 -800 175572 24
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 178966 -13 179166 46789
rect 179006 -800 179118 -13
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182508 363 182708 48594
rect 182552 -800 182664 363
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186054 326 186254 49796
rect 186098 -800 186210 326
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189594 221 189794 50868
rect 189644 -800 189756 221
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193140 11 193340 51607
rect 193190 -800 193302 11
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196697 166 196897 52370
rect 196736 -800 196848 166
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200243 129 200443 53417
rect 200282 -800 200394 129
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203783 24 203983 53882
rect 203828 -800 203940 24
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207330 -6 207530 54595
rect 207374 -800 207486 -6
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210880 363 211080 55075
rect 210920 -800 211032 363
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214426 326 214626 55599
rect 214466 -800 214578 326
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 217966 221 218166 55957
rect 218012 -800 218124 221
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221512 184 221712 56241
rect 221558 -800 221670 184
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225069 166 225269 56648
rect 225104 -800 225216 166
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228615 129 228815 57606
rect 228650 -800 228762 129
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232155 24 232355 57968
rect 232196 -800 232308 24
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235701 -13 235901 58493
rect 235742 -800 235854 -13
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239243 363 239443 61741
rect 239288 -800 239400 363
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242789 326 242989 62475
rect 242834 -800 242946 326
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246324 15 246524 63303
rect 246380 -800 246492 15
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249875 11 250075 64146
rect 249926 -800 250038 11
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253432 166 253632 65300
rect 253472 -800 253584 166
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 256978 129 257178 66596
rect 257018 -800 257130 129
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260518 24 260718 67230
rect 260564 -800 260676 24
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264065 -6 264265 69582
rect 264110 -800 264222 -6
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267615 363 267815 70469
rect 267656 -800 267768 363
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271161 326 271361 71845
rect 271202 -800 271314 326
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274701 221 274901 73190
rect 274748 -800 274860 221
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278247 184 278447 74267
rect 278294 -800 278406 184
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281804 166 282004 75085
rect 281840 -800 281952 166
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285350 129 285550 76732
rect 285386 -800 285498 129
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288890 24 289090 77783
rect 288932 -800 289044 24
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292436 -13 292636 78843
rect 292478 -800 292590 -13
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 295980 363 296180 80700
rect 296024 -800 296136 363
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299526 326 299726 82594
rect 299570 -800 299682 326
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303061 15 303261 84007
rect 303116 -800 303228 15
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306612 11 306812 84905
rect 306662 -800 306774 11
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310169 166 310369 85336
rect 310208 -800 310320 166
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313715 129 313915 85761
rect 313754 -800 313866 129
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317255 24 317455 86227
rect 317300 -800 317412 24
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320802 -6 321002 86585
rect 320846 -800 320958 -6
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324352 363 324552 86993
rect 324392 -800 324504 363
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327898 326 328098 87753
rect 327938 -800 328050 326
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331438 221 331638 88361
rect 331484 -800 331596 221
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 334984 184 335184 89004
rect 335030 -800 335142 184
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338541 166 338741 89470
rect 338576 -800 338688 166
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342087 129 342287 89756
rect 342122 -800 342234 129
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345627 24 345827 90351
rect 345668 -800 345780 24
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349173 -13 349373 91412
rect 349214 -800 349326 -13
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352705 174 352905 92796
rect 352760 -800 352872 174
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356258 174 356458 95135
rect 356306 -800 356418 174
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359801 174 360001 97918
rect 359852 -800 359964 174
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363354 174 363554 99345
rect 363398 -800 363510 174
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366892 174 367092 100482
rect 366944 -800 367056 174
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370445 174 370645 101497
rect 370490 -800 370602 174
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 373988 174 374188 102624
rect 374036 -800 374148 174
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377541 130 377741 103336
rect 381073 60383 381273 60454
rect 381073 60327 381143 60383
rect 381199 60327 381273 60383
rect 377582 -800 377694 130
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381073 174 381273 60327
rect 381128 -800 381240 174
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384626 174 384826 59357
rect 388169 58430 388369 58501
rect 388169 58374 388239 58430
rect 388295 58374 388369 58430
rect 384674 -800 384786 174
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388169 174 388369 58374
rect 391722 58027 391922 58122
rect 391722 57971 391787 58027
rect 391843 57971 391922 58027
rect 388220 -800 388332 174
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391722 174 391922 57971
rect 395260 57700 395460 57741
rect 395260 57644 395335 57700
rect 395391 57644 395460 57700
rect 391766 -800 391878 174
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395260 174 395460 57644
rect 398813 57050 399013 57080
rect 398813 56994 398880 57050
rect 398936 56994 399013 57050
rect 395312 -800 395424 174
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398813 174 399013 56994
rect 402356 56548 402556 56589
rect 402356 56492 402422 56548
rect 402478 56492 402556 56548
rect 398858 -800 398970 174
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402356 174 402556 56492
rect 405909 56033 406109 56055
rect 405909 55977 405983 56033
rect 406039 55977 406109 56033
rect 402404 -800 402516 174
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405909 174 406109 55977
rect 409458 54165 409658 54300
rect 409458 54109 409531 54165
rect 409587 54109 409658 54165
rect 405950 -800 406062 174
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409458 274 409658 54109
rect 413003 53349 413203 53505
rect 413003 53293 413076 53349
rect 413132 53293 413203 53349
rect 409496 -800 409608 274
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413003 250 413203 53293
rect 416560 52772 416760 52823
rect 416560 52716 416628 52772
rect 416684 52716 416760 52772
rect 413042 -800 413154 250
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416560 112 416760 52716
rect 420089 52250 420289 52361
rect 420089 52194 420154 52250
rect 420210 52194 420289 52250
rect 416588 -800 416700 112
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420089 271 420289 52194
rect 423643 51913 423843 52022
rect 423643 51857 423714 51913
rect 423770 51857 423843 51913
rect 420134 -800 420246 271
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423643 199 423843 51857
rect 427191 50914 427391 50975
rect 427191 50858 427266 50914
rect 427322 50858 427391 50914
rect 423680 -800 423792 199
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427191 242 427391 50858
rect 430718 50357 430918 50423
rect 430718 50301 430790 50357
rect 430846 50301 430918 50357
rect 427226 -800 427338 242
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430718 215 430918 50301
rect 434276 49414 434476 49468
rect 434276 49358 434349 49414
rect 434405 49358 434476 49414
rect 430772 -800 430884 215
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434276 223 434476 49358
rect 437809 48760 438009 48802
rect 437809 48704 437875 48760
rect 437931 48704 438009 48760
rect 434318 -800 434430 223
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437809 130 438009 48704
rect 441364 48095 441564 48171
rect 441364 48039 441438 48095
rect 441494 48039 441564 48095
rect 437864 -800 437976 130
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441364 241 441564 48039
rect 444928 47453 445128 47501
rect 444928 47397 444991 47453
rect 445047 47397 445128 47453
rect 441410 -800 441522 241
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444928 160 445128 47397
rect 448450 46925 448650 47029
rect 448450 46869 448515 46925
rect 448571 46869 448650 46925
rect 444956 -800 445068 160
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448450 152 448650 46869
rect 452010 46561 452210 46653
rect 452010 46505 452075 46561
rect 452131 46505 452210 46561
rect 448502 -800 448614 152
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452010 255 452210 46505
rect 455553 45714 455753 45765
rect 455553 45658 455623 45714
rect 455679 45658 455753 45714
rect 452048 -800 452160 255
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455553 311 455753 45658
rect 459103 45157 459303 45235
rect 459103 45101 459169 45157
rect 459225 45101 459303 45157
rect 455594 -800 455706 311
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459103 364 459303 45101
rect 462648 44462 462848 44522
rect 462648 44406 462719 44462
rect 462775 44406 462848 44462
rect 459140 -800 459252 364
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462648 199 462848 44406
rect 462686 -800 462798 199
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551291 83 551491 576269
rect 551336 -800 551448 83
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554840 84 555040 576996
rect 554882 -800 554994 84
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558390 84 558590 577586
rect 558428 -800 558540 84
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561929 159 562129 599468
rect 561974 -800 562086 159
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565471 100 565671 600723
rect 565520 -800 565632 100
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569018 200 569218 601724
rect 576111 556817 576311 571524
rect 576111 556681 576143 556817
rect 576279 556681 576311 556817
rect 572569 548905 572769 549991
rect 572569 548873 572770 548905
rect 572569 548737 572602 548873
rect 572738 548737 572770 548873
rect 572569 548705 572770 548737
rect 569066 -800 569178 200
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572569 83 572769 548705
rect 572612 -800 572724 83
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576111 201 576311 556681
rect 576158 -800 576270 201
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 538383 694684 538519 694820
rect 95449 687795 95825 687797
rect 95449 687423 95451 687795
rect 95451 687423 95823 687795
rect 95823 687423 95825 687795
rect 95449 687421 95825 687423
rect 172232 688018 172608 688020
rect 172232 687646 172234 688018
rect 172234 687646 172606 688018
rect 172606 687646 172608 688018
rect 172232 687644 172608 687646
rect 120774 687609 121150 687611
rect 120774 687237 120776 687609
rect 120776 687237 121148 687609
rect 121148 687237 121150 687609
rect 120774 687235 121150 687237
rect 146431 687487 146807 687489
rect 146431 687115 146433 687487
rect 146433 687115 146805 687487
rect 146805 687115 146807 687487
rect 146431 687113 146807 687115
rect 216370 687578 216746 687580
rect 216370 687206 216372 687578
rect 216372 687206 216744 687578
rect 216744 687206 216746 687578
rect 216370 687204 216746 687206
rect 223351 687653 223727 687655
rect 223351 687281 223353 687653
rect 223353 687281 223725 687653
rect 223725 687281 223727 687653
rect 223351 687279 223727 687281
rect 249021 687556 249397 687558
rect 249021 687184 249023 687556
rect 249023 687184 249395 687556
rect 249395 687184 249397 687556
rect 249021 687182 249397 687184
rect 274690 687572 275066 687574
rect 274690 687200 274692 687572
rect 274692 687200 275064 687572
rect 275064 687200 275066 687572
rect 274690 687198 275066 687200
rect 300315 687608 300691 687610
rect 300315 687236 300317 687608
rect 300317 687236 300689 687608
rect 300689 687236 300691 687608
rect 300315 687234 300691 687236
rect 325951 687573 326327 687575
rect 325951 687201 325953 687573
rect 325953 687201 326325 687573
rect 326325 687201 326327 687573
rect 325951 687199 326327 687201
rect 351616 687555 351992 687557
rect 351616 687183 351618 687555
rect 351618 687183 351990 687555
rect 351990 687183 351992 687555
rect 351616 687181 351992 687183
rect 377277 687517 377653 687519
rect 377277 687145 377279 687517
rect 377279 687145 377651 687517
rect 377651 687145 377653 687517
rect 377277 687143 377653 687145
rect 412453 687634 412829 687636
rect 412453 687262 412455 687634
rect 412455 687262 412827 687634
rect 412827 687262 412829 687634
rect 412453 687260 412829 687262
rect 428579 687624 428955 687626
rect 428579 687252 428581 687624
rect 428581 687252 428953 687624
rect 428953 687252 428955 687624
rect 428579 687250 428955 687252
rect 454213 687693 454589 687695
rect 454213 687321 454215 687693
rect 454215 687321 454587 687693
rect 454587 687321 454589 687693
rect 454213 687319 454589 687321
rect 479862 687699 480238 687701
rect 479862 687327 479864 687699
rect 479864 687327 480236 687699
rect 480236 687327 480238 687699
rect 479862 687325 480238 687327
rect 198548 674550 198684 674686
rect 20001 660421 20377 660797
rect 396896 660543 397032 660679
rect 416192 658802 416568 659178
rect 5039 560367 5415 560743
rect 182013 559327 182389 559703
rect 185005 559295 185381 559671
rect 186496 559304 186872 559680
rect 198430 559203 198806 559579
rect 388961 559387 389337 559763
rect 392008 559303 392384 559679
rect 393440 559289 393816 559665
rect 405364 559288 405740 559664
rect 204061 556612 204197 556748
rect 411001 556682 411137 556818
rect 24162 553247 24538 553623
rect 396896 550067 397032 550203
rect 200966 548831 201102 548967
rect 193963 548375 194099 548511
rect 37863 542331 38239 542707
rect 184194 530755 184330 530891
rect 198084 539743 198220 539879
rect 208781 539741 208917 539877
rect 201903 539235 202039 539371
rect 210004 539235 210140 539371
rect 197476 530756 197612 530892
rect 206406 530754 206542 530890
rect 391180 530756 391316 530892
rect 414690 547437 414826 547573
rect 415367 547444 415503 547580
rect 405259 539853 405395 539989
rect 408892 539401 409028 539537
rect 404425 530755 404561 530891
rect 422082 530755 422218 530891
rect 96021 445973 96157 446109
rect 76156 437887 76292 438023
rect 79804 437628 79940 437764
rect 24161 215413 24537 215789
rect 29695 225000 29831 225136
rect 273 124769 409 124905
rect 88358 435687 88494 435823
rect 80291 435488 80427 435624
rect 76173 435131 76309 435267
rect 77104 433975 77240 434111
rect 79035 433027 79171 433163
rect 76183 424547 76319 424683
rect 76198 421781 76334 421917
rect 77137 420623 77273 420759
rect 76167 411203 76303 411339
rect 76198 408436 76334 408572
rect 77125 407283 77261 407419
rect 76180 397848 76316 397984
rect 76185 395094 76321 395230
rect 77137 393934 77273 394070
rect 76155 384508 76291 384644
rect 76160 381746 76296 381882
rect 77125 380590 77261 380726
rect 76175 371166 76311 371302
rect 76178 368405 76314 368541
rect 77087 367245 77223 367381
rect 76165 357817 76301 357953
rect 76185 355060 76321 355196
rect 77177 353901 77313 354037
rect 76132 344472 76268 344608
rect 76155 341710 76291 341846
rect 79026 419680 79162 419816
rect 79010 406335 79146 406471
rect 79035 392995 79171 393131
rect 79001 379648 79137 379784
rect 79020 366299 79156 366435
rect 77143 340559 77279 340695
rect 76175 331128 76311 331264
rect 76179 328370 76315 328506
rect 77131 327216 77267 327352
rect 76187 317776 76323 317912
rect 76175 315025 76311 315161
rect 79024 352959 79160 353095
rect 79031 339610 79167 339746
rect 77136 313870 77272 314006
rect 76170 304435 76306 304571
rect 76185 301678 76321 301814
rect 77142 300519 77278 300655
rect 76170 291095 76306 291231
rect 76160 288342 76296 288478
rect 77139 287176 77275 287312
rect 76178 277761 76314 277897
rect 76178 274983 76314 275119
rect 77150 273832 77286 273968
rect 76189 264404 76325 264540
rect 76201 261645 76337 261781
rect 77152 260487 77288 260623
rect 76186 251055 76322 251191
rect 76184 248296 76320 248432
rect 77130 247140 77266 247276
rect 76233 237682 76369 237818
rect 76231 234914 76367 235050
rect 77108 233758 77244 233894
rect 76613 216167 76989 216543
rect 79043 326262 79179 326398
rect 79002 312924 79138 313060
rect 79015 299573 79151 299709
rect 79013 286230 79149 286366
rect 79020 272891 79156 273027
rect 79007 259540 79143 259676
rect 121339 254632 121475 254768
rect 79021 246194 79157 246330
rect 79016 232812 79152 232948
rect 77411 215410 77787 215786
rect 78422 214530 78798 214906
rect 96762 225000 96898 225136
rect 82023 216166 82399 216542
rect 82026 215411 82402 215787
rect 91822 215092 91958 215228
rect 104167 215083 104303 215219
rect 117141 215105 117277 215241
rect 129476 215043 129612 215179
rect 142791 215059 142927 215195
rect 155131 215089 155267 215225
rect 168433 215046 168569 215182
rect 180787 215077 180923 215213
rect 194076 215105 194212 215241
rect 206434 215083 206570 215219
rect 219731 215082 219867 215218
rect 232078 215117 232214 215253
rect 245382 215101 245518 215237
rect 257727 215132 257863 215268
rect 271036 215113 271172 215249
rect 283379 215095 283515 215231
rect 296682 215091 296818 215227
rect 309026 215098 309162 215234
rect 322333 215075 322469 215211
rect 334677 215105 334813 215241
rect 347983 215075 348119 215211
rect 360327 215087 360463 215223
rect 373632 215079 373768 215215
rect 385977 215106 386113 215242
rect 399282 215105 399418 215241
rect 411631 215071 411767 215207
rect 424931 215074 425067 215210
rect 437279 215092 437415 215228
rect 450575 215092 450711 215228
rect 462926 215079 463062 215215
rect 476238 215067 476374 215203
rect 488579 215085 488715 215221
rect 82044 214529 82420 214905
rect 79444 213740 79820 214116
rect 82058 213741 82434 214117
rect 90875 213287 91011 213423
rect 103225 213285 103361 213421
rect 116185 213286 116321 213422
rect 128528 213245 128664 213381
rect 141833 213205 141969 213341
rect 154177 213270 154313 213406
rect 167488 213231 167624 213367
rect 179832 213265 179968 213401
rect 193142 213257 193278 213393
rect 205478 213271 205614 213407
rect 218783 213272 218919 213408
rect 231133 213259 231269 213395
rect 244432 213249 244568 213385
rect 256781 213269 256917 213405
rect 270090 213250 270226 213386
rect 282434 213227 282570 213363
rect 295737 213242 295873 213378
rect 308085 213200 308221 213336
rect 321383 213259 321519 213395
rect 333728 213216 333864 213352
rect 347034 213283 347170 213419
rect 359383 213271 359519 213407
rect 372686 213283 372822 213419
rect 385033 213284 385169 213420
rect 398330 213279 398466 213415
rect 410678 213279 410814 213415
rect 423987 213282 424123 213418
rect 436212 213529 436588 213531
rect 436212 213157 436214 213529
rect 436214 213157 436586 213529
rect 436586 213157 436588 213529
rect 436212 213155 436588 213157
rect 449637 213275 449773 213411
rect 461985 213273 462121 213409
rect 475282 213268 475418 213404
rect 487630 213242 487766 213378
rect 86961 212626 87097 212762
rect 89723 212595 89859 212731
rect 99306 212575 99442 212711
rect 102079 212600 102215 212736
rect 112266 212610 112402 212746
rect 115033 212635 115169 212771
rect 124605 212600 124741 212736
rect 127378 212591 127514 212727
rect 137921 212587 138057 212723
rect 140683 212607 140819 212743
rect 150263 212548 150399 212684
rect 153021 212564 153157 212700
rect 163563 212565 163699 212701
rect 166334 212553 166470 212689
rect 175913 212572 176049 212708
rect 178674 212553 178810 212689
rect 189217 212579 189353 212715
rect 191984 212579 192120 212715
rect 201558 212589 201694 212725
rect 204324 212567 204460 212703
rect 214866 212609 215002 212745
rect 217630 212605 217766 212741
rect 227217 212598 227353 212734
rect 229976 212576 230112 212712
rect 240518 212597 240654 212733
rect 243279 212606 243415 212742
rect 252864 212587 253000 212723
rect 255624 212587 255760 212723
rect 266165 212503 266301 212639
rect 268932 212537 269068 212673
rect 278509 212568 278645 212704
rect 281277 212578 281413 212714
rect 291817 212512 291953 212648
rect 294580 212533 294716 212669
rect 304169 212553 304305 212689
rect 306933 212548 307069 212684
rect 317472 212568 317608 212704
rect 320230 212568 320366 212704
rect 329813 212595 329949 212731
rect 332576 212630 332712 212766
rect 343119 212566 343255 212702
rect 345881 212571 346017 212707
rect 355460 212562 355596 212698
rect 358226 212581 358362 212717
rect 368769 212548 368905 212684
rect 371531 212572 371667 212708
rect 381113 212595 381249 212731
rect 383878 212614 384014 212750
rect 394420 212559 394556 212695
rect 397181 212609 397317 212745
rect 406759 212575 406895 212711
rect 409528 212595 409664 212731
rect 420069 212600 420205 212736
rect 422832 212618 422968 212754
rect 432418 212615 432554 212751
rect 435177 212587 435313 212723
rect 445713 212532 445849 212668
rect 448481 212586 448617 212722
rect 458063 212547 458199 212683
rect 460825 212579 460961 212715
rect 471360 212501 471496 212637
rect 474132 212555 474268 212691
rect 483716 212513 483852 212649
rect 486479 212583 486615 212719
rect 101222 212272 101278 212328
rect 126535 212259 126591 212315
rect 100258 192038 100314 192094
rect 125563 191875 125619 191931
rect 152186 212258 152242 212314
rect 151219 189899 151275 189955
rect 177825 212254 177881 212310
rect 176862 190269 176918 190325
rect 203481 212260 203537 212316
rect 202501 188057 202557 188113
rect 229120 212260 229176 212316
rect 228168 187350 228224 187406
rect 254787 212257 254843 212313
rect 253806 188659 253862 188715
rect 280430 212260 280486 212316
rect 279460 186881 279516 186937
rect 306083 212255 306139 212311
rect 305111 186316 305167 186372
rect 331729 212255 331785 212311
rect 330761 187353 330817 187409
rect 357376 212264 357432 212320
rect 356415 189596 356471 189652
rect 383011 212260 383067 212316
rect 382053 190974 382109 191030
rect 408677 212260 408733 212316
rect 407725 192321 407781 192377
rect 434314 212255 434370 212311
rect 433370 194455 433426 194511
rect 459979 212256 460035 212312
rect 459011 195870 459067 195926
rect 485620 212258 485676 212314
rect 484658 197044 484714 197100
rect 377607 103336 377663 103392
rect 374062 102624 374118 102680
rect 370515 101497 370571 101553
rect 366968 100482 367024 100538
rect 363423 99345 363479 99401
rect 359877 97918 359933 97974
rect 356344 95135 356400 95191
rect 352774 92796 352830 92852
rect 381143 60327 381199 60383
rect 388239 58374 388295 58430
rect 391787 57971 391843 58027
rect 395335 57644 395391 57700
rect 398880 56994 398936 57050
rect 402422 56492 402478 56548
rect 405983 55977 406039 56033
rect 409531 54109 409587 54165
rect 413076 53293 413132 53349
rect 416628 52716 416684 52772
rect 420154 52194 420210 52250
rect 423714 51857 423770 51913
rect 427266 50858 427322 50914
rect 430790 50301 430846 50357
rect 434349 49358 434405 49414
rect 437875 48704 437931 48760
rect 441438 48039 441494 48095
rect 444991 47397 445047 47453
rect 448515 46869 448571 46925
rect 452075 46505 452131 46561
rect 455623 45658 455679 45714
rect 459169 45101 459225 45157
rect 462719 44406 462775 44462
rect 576143 556681 576279 556817
rect 572602 548737 572738 548873
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 18937 697229 19337 702300
rect 18937 696829 61485 697229
rect -800 683156 1700 685242
rect -800 682756 20377 683156
rect -800 680242 1700 682756
rect 19977 660809 20377 682756
rect 61085 671400 61485 696829
rect 70354 674457 70754 702300
rect 95437 687801 95837 687809
rect 95437 687417 95445 687801
rect 95829 687417 95837 687801
rect 95437 687409 95837 687417
rect 120762 687615 121162 687623
rect 120762 687231 120770 687615
rect 121154 687231 121162 687615
rect 120762 687223 121162 687231
rect 122342 676466 122742 702300
rect 167706 699875 168106 702300
rect 171703 699875 172103 699877
rect 178185 699875 178585 702300
rect 167706 699475 178585 699875
rect 219242 699612 219642 702300
rect 223956 699612 224356 699614
rect 230371 699612 230771 702300
rect 146419 687493 146819 687501
rect 146419 687109 146427 687493
rect 146811 687109 146819 687493
rect 146419 687101 146819 687109
rect 171703 681551 172103 699475
rect 219242 699212 230771 699612
rect 223956 691375 224356 699212
rect 321036 697404 321436 702300
rect 332256 697404 332656 702300
rect 321036 697004 332656 697404
rect 223956 690975 265668 691375
rect 172220 688024 172620 688032
rect 172220 687640 172228 688024
rect 172612 687640 172620 688024
rect 172220 687632 172620 687640
rect 223339 687659 223739 687667
rect 216358 687584 216758 687592
rect 216358 687200 216366 687584
rect 216750 687200 216758 687584
rect 223339 687275 223347 687659
rect 223731 687275 223739 687659
rect 223339 687267 223739 687275
rect 249009 687562 249409 687570
rect 216358 687192 216758 687200
rect 249009 687178 249017 687562
rect 249401 687178 249409 687562
rect 249009 687170 249409 687178
rect 171703 681151 255445 681551
rect 122342 676066 186871 676466
rect 70354 674057 185387 674457
rect 61085 671000 182398 671400
rect 19977 660797 20389 660809
rect 19977 660421 20001 660797
rect 20377 660421 20389 660797
rect 19977 660409 20389 660421
rect 19977 660315 20377 660409
rect -800 646503 1660 648642
rect -800 646103 24549 646503
rect -800 643842 1660 646103
rect -800 633842 1660 638642
rect -800 560757 1660 564242
rect -800 560743 5431 560757
rect -800 560367 5039 560743
rect 5415 560367 5431 560743
rect -800 560357 5431 560367
rect -800 559442 1660 560357
rect 5027 560355 5427 560357
rect -800 549442 1660 554242
rect 24149 553635 24549 646103
rect 181998 559715 182398 671000
rect 181998 559703 182401 559715
rect 181998 559327 182013 559703
rect 182389 559327 182401 559703
rect 181998 559315 182401 559327
rect 184987 559683 185387 674057
rect 186471 559692 186871 676066
rect 198419 674686 198819 674822
rect 198419 674550 198548 674686
rect 198684 674550 198819 674686
rect 184987 559671 185393 559683
rect 181998 559312 182398 559315
rect 184987 559295 185005 559671
rect 185381 559295 185393 559671
rect 184987 559288 185393 559295
rect 186471 559680 186884 559692
rect 186471 559304 186496 559680
rect 186872 559304 186884 559680
rect 198419 559591 198819 674550
rect 255045 575066 255445 681151
rect 265268 577745 265668 690975
rect 300303 687614 300703 687622
rect 274678 687578 275078 687586
rect 274678 687194 274686 687578
rect 275070 687194 275078 687578
rect 300303 687230 300311 687614
rect 300695 687230 300703 687614
rect 300303 687222 300703 687230
rect 274678 687186 275078 687194
rect 322770 592312 323170 697004
rect 412441 687640 412841 687648
rect 325939 687579 326339 687587
rect 325939 687195 325947 687579
rect 326331 687195 326339 687579
rect 325939 687187 326339 687195
rect 351604 687561 352004 687569
rect 351604 687177 351612 687561
rect 351996 687177 352004 687561
rect 351604 687169 352004 687177
rect 377265 687523 377665 687531
rect 377265 687139 377273 687523
rect 377657 687139 377665 687523
rect 412441 687256 412449 687640
rect 412833 687256 412841 687640
rect 412441 687248 412841 687256
rect 377265 687131 377665 687139
rect 396864 660679 397064 660807
rect 396864 660543 396896 660679
rect 397032 660543 397064 660679
rect 322770 591912 393804 592312
rect 265268 577345 392377 577745
rect 255045 574666 389355 575066
rect 388955 559775 389355 574666
rect 186471 559292 186884 559304
rect 198418 559579 198819 559591
rect 186471 559291 186871 559292
rect 184993 559283 185393 559288
rect 198418 559203 198430 559579
rect 198806 559203 198819 559579
rect 388949 559763 389355 559775
rect 388949 559387 388961 559763
rect 389337 559387 389355 559763
rect 388949 559375 389355 559387
rect 388955 559372 389355 559375
rect 391977 559691 392377 577345
rect 391977 559679 392396 559691
rect 198418 559191 198819 559203
rect 391977 559303 392008 559679
rect 392384 559303 392396 559679
rect 391977 559291 392396 559303
rect 393404 559677 393804 591912
rect 393404 559665 393828 559677
rect 391977 559194 392377 559291
rect 393404 559289 393440 559665
rect 393816 559289 393828 559665
rect 393404 559277 393828 559289
rect 198419 559190 198819 559191
rect 393404 559185 393804 559277
rect 203992 556748 214191 556780
rect 203992 556612 204061 556748
rect 204197 556612 214191 556748
rect 203992 556580 214191 556612
rect 24149 553623 24550 553635
rect 24149 553247 24162 553623
rect 24538 553247 24550 553623
rect 24149 553235 24550 553247
rect 24149 553233 24549 553235
rect 6084 548967 201149 548999
rect 6084 548831 200966 548967
rect 201102 548831 201149 548967
rect 6084 548799 201149 548831
rect 213991 548904 214191 556580
rect 396864 550203 397064 660543
rect 416179 659190 416579 702300
rect 510594 688454 515394 704800
rect 454201 687699 454601 687707
rect 428567 687630 428967 687638
rect 428567 687246 428575 687630
rect 428959 687246 428967 687630
rect 454201 687315 454209 687699
rect 454593 687315 454601 687699
rect 454201 687307 454601 687315
rect 479850 687705 480250 687713
rect 479850 687321 479858 687705
rect 480242 687321 480250 687705
rect 479850 687313 480250 687321
rect 510594 687670 512525 688454
rect 513309 687670 515394 688454
rect 428567 687238 428967 687246
rect 416179 659178 416580 659190
rect 416179 658802 416192 659178
rect 416568 658802 416580 659178
rect 416179 658790 416580 658802
rect 510594 631116 515394 687670
rect 520594 688496 525394 704800
rect 566594 702300 571594 704800
rect 568970 694957 569370 702300
rect 538246 694820 569370 694957
rect 538246 694684 538383 694820
rect 538519 694684 569370 694820
rect 538246 694557 569370 694684
rect 520594 687712 522690 688496
rect 523474 687712 525394 688496
rect 520594 631116 525394 687712
rect 582300 680616 584800 682984
rect 544336 680216 584800 680616
rect 544336 559676 544736 680216
rect 582300 677984 584800 680216
rect 560050 644576 584800 644584
rect 560050 639792 560582 644576
rect 566726 639792 584800 644576
rect 560050 639784 584800 639792
rect 560050 634576 584800 634584
rect 560050 629792 560582 634576
rect 566726 629792 584800 634576
rect 560050 629784 584800 629792
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 405314 559664 544736 559676
rect 405314 559288 405364 559664
rect 405740 559288 544736 559664
rect 405314 559276 544736 559288
rect 410938 556818 576311 556850
rect 410938 556682 411001 556818
rect 411137 556817 576311 556818
rect 411137 556682 576143 556817
rect 410938 556681 576143 556682
rect 576279 556681 576311 556817
rect 410938 556650 576311 556681
rect 576111 556649 576311 556650
rect 555452 555354 584800 555362
rect 555452 550570 556255 555354
rect 562319 550570 584800 555354
rect 555452 550562 584800 550570
rect 396864 550067 396896 550203
rect 397032 550067 397064 550203
rect 396864 549891 397064 550067
rect 572570 548904 572770 548905
rect 213991 548873 572773 548904
rect 6084 511683 6284 548799
rect 213991 548737 572602 548873
rect 572738 548737 572773 548873
rect 213991 548704 572773 548737
rect 466 511642 6284 511683
rect -800 511530 6284 511642
rect 466 511483 6284 511530
rect 6965 548543 194087 548544
rect 6965 548511 194131 548543
rect 6965 548375 193963 548511
rect 194099 548375 194131 548511
rect 6965 548344 194131 548375
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 6965 468447 7165 548344
rect 193931 548343 194131 548344
rect 414658 547573 414858 547656
rect 414658 547437 414690 547573
rect 414826 547437 414858 547573
rect 37851 542711 38251 542719
rect 37851 542327 37859 542711
rect 38243 542327 38251 542711
rect 37851 542319 38251 542327
rect 414658 540021 414858 547437
rect 404978 539989 414858 540021
rect 197943 539879 209042 539911
rect 197943 539743 198084 539879
rect 198220 539877 209042 539879
rect 198220 539743 208781 539877
rect 197943 539741 208781 539743
rect 208917 539741 209042 539877
rect 404978 539853 405259 539989
rect 405395 539853 414858 539989
rect 404978 539821 414858 539853
rect 415335 547580 415535 547660
rect 415335 547444 415367 547580
rect 415503 547444 415535 547580
rect 197943 539711 209042 539741
rect 208749 539709 208949 539711
rect 415335 539569 415535 547444
rect 555452 545354 584800 545362
rect 555452 540570 556255 545354
rect 562319 540570 584800 545354
rect 555452 540562 584800 540570
rect 408739 539537 415535 539569
rect 201773 539371 210360 539403
rect 201773 539235 201903 539371
rect 202039 539235 210004 539371
rect 210140 539235 210360 539371
rect 408739 539401 408892 539537
rect 409028 539401 415535 539537
rect 408739 539369 415535 539401
rect 201773 539203 210360 539235
rect 10426 531016 10826 531024
rect 10426 530923 10434 531016
rect 9941 530723 10434 530923
rect 10426 530632 10434 530723
rect 10818 530923 10826 531016
rect 569780 531017 570180 531025
rect 197444 530923 197644 530924
rect 391148 530923 391348 530924
rect 569780 530923 569788 531017
rect 10818 530892 569788 530923
rect 10818 530891 197476 530892
rect 10818 530755 184194 530891
rect 184330 530756 197476 530891
rect 197612 530890 391180 530892
rect 197612 530756 206406 530890
rect 184330 530755 206406 530756
rect 10818 530754 206406 530755
rect 206542 530756 391180 530890
rect 391316 530891 569788 530892
rect 391316 530756 404425 530891
rect 206542 530755 404425 530756
rect 404561 530755 422082 530891
rect 422218 530755 569788 530891
rect 206542 530754 569788 530755
rect 10818 530723 569788 530754
rect 10818 530632 10826 530723
rect 206374 530722 206574 530723
rect 10426 530624 10826 530632
rect 569780 530633 569788 530723
rect 570172 530923 570180 531017
rect 570172 530723 570387 530923
rect 570172 530633 570180 530723
rect 569780 530625 570180 530633
rect 573371 500050 583220 500162
rect 583318 500050 584800 500162
rect 539494 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 410 468420 7165 468447
rect -800 468308 7165 468420
rect 410 468247 7165 468308
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 660 462510
rect 780 462398 17711 462510
rect 573405 455628 583180 455740
rect 583296 455628 584800 455740
rect 537376 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 3838 446109 96189 446142
rect 3838 445973 96021 446109
rect 96157 445973 96189 446109
rect 3838 445942 96189 445973
rect 3838 425244 4038 445942
rect 95989 445941 96189 445942
rect 393 425198 4038 425244
rect -800 425086 4038 425198
rect 393 425044 4038 425086
rect 20602 444360 88525 444560
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 676 419288
rect 738 419176 17694 419288
rect 20602 382035 20802 444360
rect 352 381976 20802 382035
rect -800 381864 20802 381976
rect 352 381835 20802 381864
rect 22298 442803 80459 443003
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 22298 338784 22498 442803
rect 287 338754 22498 338784
rect -800 338642 22498 338754
rect 287 338584 22498 338642
rect 26220 440887 79971 441087
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 26220 295556 26420 440887
rect 76124 438027 76324 438055
rect 76124 437883 76152 438027
rect 76296 437883 76324 438027
rect 76124 437855 76324 437883
rect 79771 437796 79971 440887
rect 79771 437764 79972 437796
rect 79771 437628 79804 437764
rect 79940 437628 79972 437764
rect 79771 437597 79972 437628
rect 79772 437596 79972 437597
rect 80259 435624 80459 442803
rect 88325 435855 88525 444360
rect 88325 435823 88526 435855
rect 88325 435687 88358 435823
rect 88494 435687 88526 435823
rect 88325 435655 88526 435687
rect 88325 435635 88525 435655
rect 80259 435488 80291 435624
rect 80427 435488 80459 435624
rect 80259 435456 80459 435488
rect 76141 435271 76341 435299
rect 76141 435127 76169 435271
rect 76313 435127 76341 435271
rect 76141 435099 76341 435127
rect 77072 434115 77272 434143
rect 77072 433971 77100 434115
rect 77244 433971 77272 434115
rect 77072 433943 77272 433971
rect 79003 433167 79203 433195
rect 79003 433023 79031 433167
rect 79175 433023 79203 433167
rect 79003 432995 79203 433023
rect 76151 424687 76351 424715
rect 76151 424543 76179 424687
rect 76323 424543 76351 424687
rect 76151 424515 76351 424543
rect 76166 421921 76366 421949
rect 76166 421777 76194 421921
rect 76338 421777 76366 421921
rect 76166 421749 76366 421777
rect 77105 420763 77305 420791
rect 77105 420619 77133 420763
rect 77277 420619 77305 420763
rect 77105 420591 77305 420619
rect 78994 419820 79194 419848
rect 78994 419676 79022 419820
rect 79166 419676 79194 419820
rect 78994 419648 79194 419676
rect 76135 411343 76335 411371
rect 76135 411199 76163 411343
rect 76307 411199 76335 411343
rect 583520 411206 584800 411318
rect 76135 411171 76335 411199
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 76166 408576 76366 408604
rect 76166 408432 76194 408576
rect 76338 408432 76366 408576
rect 76166 408404 76366 408432
rect 583520 407660 584800 407772
rect 77093 407423 77293 407451
rect 77093 407279 77121 407423
rect 77265 407279 77293 407423
rect 77093 407251 77293 407279
rect 78978 406475 79178 406503
rect 583520 406478 584800 406590
rect 78978 406331 79006 406475
rect 79150 406331 79178 406475
rect 78978 406303 79178 406331
rect 533497 405296 584800 405408
rect 76148 397988 76348 398016
rect 76148 397844 76176 397988
rect 76320 397844 76348 397988
rect 76148 397816 76348 397844
rect 76153 395234 76353 395262
rect 76153 395090 76181 395234
rect 76325 395090 76353 395234
rect 76153 395062 76353 395090
rect 77105 394074 77305 394102
rect 77105 393930 77133 394074
rect 77277 393930 77305 394074
rect 77105 393902 77305 393930
rect 79003 393135 79203 393163
rect 79003 392991 79031 393135
rect 79175 392991 79203 393135
rect 79003 392963 79203 392991
rect 76123 384648 76323 384676
rect 76123 384504 76151 384648
rect 76295 384504 76323 384648
rect 76123 384476 76323 384504
rect 76128 381886 76328 381914
rect 76128 381742 76156 381886
rect 76300 381742 76328 381886
rect 76128 381714 76328 381742
rect 77093 380730 77293 380758
rect 77093 380586 77121 380730
rect 77265 380586 77293 380730
rect 77093 380558 77293 380586
rect 78969 379788 79169 379816
rect 78969 379644 78997 379788
rect 79141 379644 79169 379788
rect 78969 379616 79169 379644
rect 76143 371306 76343 371334
rect 76143 371162 76171 371306
rect 76315 371162 76343 371306
rect 76143 371134 76343 371162
rect 76146 368545 76346 368573
rect 76146 368401 76174 368545
rect 76318 368401 76346 368545
rect 76146 368373 76346 368401
rect 77055 367385 77255 367413
rect 77055 367241 77083 367385
rect 77227 367241 77255 367385
rect 77055 367213 77255 367241
rect 78988 366439 79188 366467
rect 78988 366295 79016 366439
rect 79160 366295 79188 366439
rect 78988 366267 79188 366295
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 76133 357957 76333 357985
rect 76133 357813 76161 357957
rect 76305 357813 76333 357957
rect 76133 357785 76333 357813
rect 76153 355200 76353 355228
rect 76153 355056 76181 355200
rect 76325 355056 76353 355200
rect 76153 355028 76353 355056
rect 77145 354041 77345 354069
rect 77145 353897 77173 354041
rect 77317 353897 77345 354041
rect 77145 353869 77345 353897
rect 78992 353099 79192 353127
rect 78992 352955 79020 353099
rect 79164 352955 79192 353099
rect 78992 352927 79192 352955
rect 76100 344612 76300 344640
rect 76100 344468 76128 344612
rect 76272 344468 76300 344612
rect 76100 344440 76300 344468
rect 76123 341850 76323 341878
rect 76123 341706 76151 341850
rect 76295 341706 76323 341850
rect 76123 341678 76323 341706
rect 77111 340699 77311 340727
rect 77111 340555 77139 340699
rect 77283 340555 77311 340699
rect 77111 340527 77311 340555
rect 78999 339750 79199 339778
rect 78999 339606 79027 339750
rect 79171 339606 79199 339750
rect 78999 339578 79199 339606
rect 76143 331268 76343 331296
rect 76143 331124 76171 331268
rect 76315 331124 76343 331268
rect 76143 331096 76343 331124
rect 76147 328510 76347 328538
rect 76147 328366 76175 328510
rect 76319 328366 76347 328510
rect 76147 328338 76347 328366
rect 77099 327356 77299 327384
rect 77099 327212 77127 327356
rect 77271 327212 77299 327356
rect 77099 327184 77299 327212
rect 79011 326402 79211 326430
rect 79011 326258 79039 326402
rect 79183 326258 79211 326402
rect 79011 326230 79211 326258
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 76155 317916 76355 317944
rect 76155 317772 76183 317916
rect 76327 317772 76355 317916
rect 76155 317744 76355 317772
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 76143 315165 76343 315193
rect 76143 315021 76171 315165
rect 76315 315021 76343 315165
rect 76143 314993 76343 315021
rect 583520 314834 584800 314946
rect 77104 314010 77304 314038
rect 77104 313866 77132 314010
rect 77276 313866 77304 314010
rect 77104 313838 77304 313866
rect 583520 313652 584800 313764
rect 78970 313064 79170 313092
rect 78970 312920 78998 313064
rect 79142 312920 79170 313064
rect 78970 312892 79170 312920
rect 76138 304575 76338 304603
rect 76138 304431 76166 304575
rect 76310 304431 76338 304575
rect 76138 304403 76338 304431
rect 76153 301818 76353 301846
rect 76153 301674 76181 301818
rect 76325 301674 76353 301818
rect 76153 301646 76353 301674
rect 77110 300659 77310 300687
rect 77110 300515 77138 300659
rect 77282 300515 77310 300659
rect 77110 300487 77310 300515
rect 78983 299713 79183 299741
rect 78983 299569 79011 299713
rect 79155 299569 79183 299713
rect 78983 299541 79183 299569
rect 203 295532 26420 295556
rect -800 295420 26420 295532
rect 203 295356 26420 295420
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect 76138 291235 76338 291263
rect 76138 291091 76166 291235
rect 76310 291091 76338 291235
rect 76138 291063 76338 291091
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 76128 288482 76328 288510
rect 76128 288338 76156 288482
rect 76300 288338 76328 288482
rect 76128 288310 76328 288338
rect 77107 287316 77307 287344
rect 77107 287172 77135 287316
rect 77279 287172 77307 287316
rect 77107 287144 77307 287172
rect 78981 286370 79181 286398
rect 78981 286226 79009 286370
rect 79153 286226 79181 286370
rect 78981 286198 79181 286226
rect 76146 277901 76346 277929
rect 76146 277757 76174 277901
rect 76318 277757 76346 277901
rect 76146 277729 76346 277757
rect 76146 275123 76346 275151
rect 583520 275140 584800 275252
rect 76146 274979 76174 275123
rect 76318 274979 76346 275123
rect 76146 274951 76346 274979
rect 77118 273972 77318 274000
rect 77118 273828 77146 273972
rect 77290 273828 77318 273972
rect 583520 273958 584800 274070
rect 77118 273800 77318 273828
rect 78988 273031 79188 273059
rect 78988 272887 79016 273031
rect 79160 272887 79188 273031
rect 78988 272859 79188 272887
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 76157 264544 76357 264572
rect 76157 264400 76185 264544
rect 76329 264400 76357 264544
rect 76157 264372 76357 264400
rect 76169 261785 76369 261813
rect 76169 261641 76197 261785
rect 76341 261641 76369 261785
rect 76169 261613 76369 261641
rect 77120 260627 77320 260655
rect 77120 260483 77148 260627
rect 77292 260483 77320 260627
rect 77120 260455 77320 260483
rect 78975 259680 79175 259708
rect 78975 259536 79003 259680
rect 79147 259536 79175 259680
rect 78975 259508 79175 259536
rect 1167 254768 121508 254800
rect 1167 254632 121339 254768
rect 121475 254632 121508 254768
rect 1167 254600 121508 254632
rect 1167 252553 1367 254600
rect 338 252510 1367 252553
rect -800 252398 1367 252510
rect 338 252353 1367 252398
rect -800 251216 480 251328
rect 76154 251195 76354 251223
rect 76154 251051 76182 251195
rect 76326 251051 76354 251195
rect 76154 251023 76354 251051
rect -800 250034 480 250146
rect -800 248852 480 248964
rect 76152 248436 76352 248464
rect 76152 248292 76180 248436
rect 76324 248292 76352 248436
rect 76152 248264 76352 248292
rect -800 247670 480 247782
rect 77098 247280 77298 247308
rect 77098 247136 77126 247280
rect 77270 247136 77298 247280
rect 77098 247108 77298 247136
rect -800 246488 480 246600
rect 78989 246334 79189 246362
rect 78989 246190 79017 246334
rect 79161 246190 79189 246334
rect 78989 246162 79189 246190
rect 582340 238072 584800 240030
rect 76201 237822 76401 237850
rect 76201 237678 76229 237822
rect 76373 237678 76401 237822
rect 76201 237650 76401 237678
rect 578979 237272 584800 238072
rect 76199 235054 76399 235082
rect 76199 234910 76227 235054
rect 76371 234910 76399 235054
rect 76199 234882 76399 234910
rect 77076 233898 77276 233926
rect 77076 233754 77104 233898
rect 77248 233754 77276 233898
rect 77076 233726 77276 233754
rect 578979 233680 579779 237272
rect 582340 235230 584800 237272
rect 538783 233284 579779 233680
rect 78984 232952 79184 232980
rect 78984 232808 79012 232952
rect 79156 232808 79184 232952
rect 78984 232780 79184 232808
rect 538783 231700 539194 233284
rect 540778 231700 579779 233284
rect 538783 231280 579779 231700
rect 578979 227650 579779 231280
rect 582340 227650 584800 230030
rect 578979 226850 584800 227650
rect 582340 225230 584800 226850
rect 29600 225136 96930 225169
rect 29600 225000 29695 225136
rect 29831 225000 96762 225136
rect 96898 225000 96930 225136
rect 29600 224969 96930 225000
rect 29663 224968 29863 224969
rect 96730 224968 96930 224969
rect -800 216556 1660 219688
rect -800 216543 82453 216556
rect -800 216167 76613 216543
rect 76989 216542 82453 216543
rect 76989 216167 82023 216542
rect -800 216166 82023 216167
rect 82399 216166 82453 216542
rect -800 216156 82453 216166
rect -800 214888 1660 216156
rect -800 207780 1660 209688
rect 3209 207780 3609 216156
rect 76601 216155 77001 216156
rect 82011 216154 82411 216156
rect 24149 215799 24549 215801
rect 24149 215789 82424 215799
rect 24149 215413 24161 215789
rect 24537 215787 82424 215789
rect 24537 215786 82026 215787
rect 24537 215413 77411 215786
rect 24149 215410 77411 215413
rect 77787 215411 82026 215786
rect 82402 215411 82424 215787
rect 77787 215410 82424 215411
rect 24149 215401 82424 215410
rect 24159 215399 82424 215401
rect 77399 215398 77799 215399
rect 91790 215232 91990 215260
rect 91790 215088 91818 215232
rect 91962 215088 91990 215232
rect 91790 215060 91990 215088
rect 104135 215223 104335 215251
rect 104135 215079 104163 215223
rect 104307 215079 104335 215223
rect 104135 215051 104335 215079
rect 117109 215245 117309 215273
rect 117109 215101 117137 215245
rect 117281 215101 117309 215245
rect 155099 215229 155299 215257
rect 194044 215245 194244 215273
rect 232046 215257 232246 215285
rect 257695 215272 257895 215300
rect 117109 215073 117309 215101
rect 129444 215183 129644 215211
rect 129444 215039 129472 215183
rect 129616 215039 129644 215183
rect 129444 215011 129644 215039
rect 142759 215199 142959 215227
rect 142759 215055 142787 215199
rect 142931 215055 142959 215199
rect 155099 215085 155127 215229
rect 155271 215085 155299 215229
rect 180755 215217 180955 215245
rect 155099 215057 155299 215085
rect 168401 215186 168601 215214
rect 142759 215027 142959 215055
rect 168401 215042 168429 215186
rect 168573 215042 168601 215186
rect 180755 215073 180783 215217
rect 180927 215073 180955 215217
rect 194044 215101 194072 215245
rect 194216 215101 194244 215245
rect 194044 215073 194244 215101
rect 206402 215223 206602 215251
rect 206402 215079 206430 215223
rect 206574 215079 206602 215223
rect 180755 215045 180955 215073
rect 206402 215051 206602 215079
rect 219699 215222 219899 215250
rect 219699 215078 219727 215222
rect 219871 215078 219899 215222
rect 232046 215113 232074 215257
rect 232218 215113 232246 215257
rect 232046 215085 232246 215113
rect 245350 215241 245550 215269
rect 245350 215097 245378 215241
rect 245522 215097 245550 215241
rect 257695 215128 257723 215272
rect 257867 215128 257895 215272
rect 257695 215100 257895 215128
rect 271004 215253 271204 215281
rect 271004 215109 271032 215253
rect 271176 215109 271204 215253
rect 219699 215050 219899 215078
rect 245350 215069 245550 215097
rect 271004 215081 271204 215109
rect 283347 215235 283547 215263
rect 283347 215091 283375 215235
rect 283519 215091 283547 215235
rect 283347 215063 283547 215091
rect 296650 215231 296850 215259
rect 296650 215087 296678 215231
rect 296822 215087 296850 215231
rect 296650 215059 296850 215087
rect 308994 215238 309194 215266
rect 334645 215245 334845 215273
rect 308994 215094 309022 215238
rect 309166 215094 309194 215238
rect 308994 215066 309194 215094
rect 322301 215215 322501 215243
rect 322301 215071 322329 215215
rect 322473 215071 322501 215215
rect 334645 215101 334673 215245
rect 334817 215101 334845 215245
rect 334645 215073 334845 215101
rect 347951 215215 348151 215243
rect 322301 215043 322501 215071
rect 347951 215071 347979 215215
rect 348123 215071 348151 215215
rect 347951 215043 348151 215071
rect 360295 215227 360495 215255
rect 360295 215083 360323 215227
rect 360467 215083 360495 215227
rect 360295 215055 360495 215083
rect 373600 215219 373800 215247
rect 373600 215075 373628 215219
rect 373772 215075 373800 215219
rect 373600 215047 373800 215075
rect 385945 215246 386145 215274
rect 385945 215102 385973 215246
rect 386117 215102 386145 215246
rect 385945 215074 386145 215102
rect 399250 215245 399450 215273
rect 399250 215101 399278 215245
rect 399422 215101 399450 215245
rect 399250 215073 399450 215101
rect 411599 215211 411799 215239
rect 411599 215067 411627 215211
rect 411771 215067 411799 215211
rect 168401 215014 168601 215042
rect 411599 215039 411799 215067
rect 424899 215214 425099 215242
rect 424899 215070 424927 215214
rect 425071 215070 425099 215214
rect 424899 215042 425099 215070
rect 437247 215232 437447 215260
rect 437247 215088 437275 215232
rect 437419 215088 437447 215232
rect 437247 215060 437447 215088
rect 450543 215232 450743 215260
rect 450543 215088 450571 215232
rect 450715 215088 450743 215232
rect 450543 215060 450743 215088
rect 462894 215219 463094 215247
rect 462894 215075 462922 215219
rect 463066 215075 463094 215219
rect 462894 215047 463094 215075
rect 476206 215207 476406 215235
rect 476206 215063 476234 215207
rect 476378 215063 476406 215207
rect 476206 215035 476406 215063
rect 488547 215225 488747 215253
rect 488547 215081 488575 215225
rect 488719 215081 488747 215225
rect 488547 215053 488747 215081
rect 9834 214918 10234 214919
rect 8944 214911 82592 214918
rect 8944 214527 9842 214911
rect 10226 214906 82592 214911
rect 10226 214530 78422 214906
rect 78798 214905 82592 214906
rect 78798 214530 82044 214905
rect 10226 214529 82044 214530
rect 82420 214529 82592 214905
rect 10226 214527 82592 214529
rect 8944 214518 82592 214527
rect 82032 214517 82432 214518
rect 79431 214117 82556 214129
rect 79431 214116 82058 214117
rect 79431 213740 79444 214116
rect 79820 213741 82058 214116
rect 82434 213741 82556 214117
rect 79820 213740 82556 213741
rect 79431 213729 82556 213740
rect 79432 213728 79832 213729
rect 569521 213546 569921 213547
rect 436200 213535 436600 213543
rect 90843 213427 91043 213455
rect 90843 213283 90871 213427
rect 91015 213283 91043 213427
rect 90843 213255 91043 213283
rect 103193 213425 103393 213453
rect 103193 213281 103221 213425
rect 103365 213281 103393 213425
rect 103193 213253 103393 213281
rect 116153 213426 116353 213454
rect 116153 213282 116181 213426
rect 116325 213282 116353 213426
rect 116153 213254 116353 213282
rect 128496 213385 128696 213413
rect 128496 213241 128524 213385
rect 128668 213241 128696 213385
rect 154145 213410 154345 213438
rect 128496 213213 128696 213241
rect 141801 213345 142001 213373
rect 141801 213201 141829 213345
rect 141973 213201 142001 213345
rect 154145 213266 154173 213410
rect 154317 213266 154345 213410
rect 179800 213405 180000 213433
rect 154145 213238 154345 213266
rect 167456 213371 167656 213399
rect 141801 213173 142001 213201
rect 167456 213227 167484 213371
rect 167628 213227 167656 213371
rect 179800 213261 179828 213405
rect 179972 213261 180000 213405
rect 179800 213233 180000 213261
rect 193110 213397 193310 213425
rect 193110 213253 193138 213397
rect 193282 213253 193310 213397
rect 167456 213199 167656 213227
rect 193110 213225 193310 213253
rect 205446 213411 205646 213439
rect 205446 213267 205474 213411
rect 205618 213267 205646 213411
rect 205446 213239 205646 213267
rect 218751 213412 218951 213440
rect 218751 213268 218779 213412
rect 218923 213268 218951 213412
rect 218751 213240 218951 213268
rect 231101 213399 231301 213427
rect 231101 213255 231129 213399
rect 231273 213255 231301 213399
rect 231101 213227 231301 213255
rect 244400 213389 244600 213417
rect 244400 213245 244428 213389
rect 244572 213245 244600 213389
rect 244400 213217 244600 213245
rect 256749 213409 256949 213437
rect 256749 213265 256777 213409
rect 256921 213265 256949 213409
rect 256749 213237 256949 213265
rect 270058 213390 270258 213418
rect 270058 213246 270086 213390
rect 270230 213246 270258 213390
rect 270058 213218 270258 213246
rect 282402 213367 282602 213395
rect 282402 213223 282430 213367
rect 282574 213223 282602 213367
rect 282402 213195 282602 213223
rect 295705 213382 295905 213410
rect 295705 213238 295733 213382
rect 295877 213238 295905 213382
rect 321351 213399 321551 213427
rect 295705 213210 295905 213238
rect 308053 213340 308253 213368
rect 308053 213196 308081 213340
rect 308225 213196 308253 213340
rect 321351 213255 321379 213399
rect 321523 213255 321551 213399
rect 347002 213423 347202 213451
rect 321351 213227 321551 213255
rect 333696 213356 333896 213384
rect 308053 213168 308253 213196
rect 333696 213212 333724 213356
rect 333868 213212 333896 213356
rect 347002 213279 347030 213423
rect 347174 213279 347202 213423
rect 347002 213251 347202 213279
rect 359351 213411 359551 213439
rect 359351 213267 359379 213411
rect 359523 213267 359551 213411
rect 359351 213239 359551 213267
rect 372654 213423 372854 213451
rect 372654 213279 372682 213423
rect 372826 213279 372854 213423
rect 372654 213251 372854 213279
rect 385001 213424 385201 213452
rect 385001 213280 385029 213424
rect 385173 213280 385201 213424
rect 385001 213252 385201 213280
rect 398298 213419 398498 213447
rect 398298 213275 398326 213419
rect 398470 213275 398498 213419
rect 398298 213247 398498 213275
rect 410646 213419 410846 213447
rect 410646 213275 410674 213419
rect 410818 213275 410846 213419
rect 410646 213247 410846 213275
rect 423955 213422 424155 213450
rect 423955 213278 423983 213422
rect 424127 213278 424155 213422
rect 423955 213250 424155 213278
rect 333696 213184 333896 213212
rect 436200 213151 436208 213535
rect 436592 213151 436600 213535
rect 534518 213539 570645 213546
rect 534518 213538 569529 213539
rect 449605 213415 449805 213443
rect 449605 213271 449633 213415
rect 449777 213271 449805 213415
rect 449605 213243 449805 213271
rect 461953 213413 462153 213441
rect 461953 213269 461981 213413
rect 462125 213269 462153 213413
rect 461953 213241 462153 213269
rect 475250 213408 475450 213436
rect 475250 213264 475278 213408
rect 475422 213264 475450 213408
rect 475250 213236 475450 213264
rect 487598 213382 487798 213410
rect 487598 213238 487626 213382
rect 487770 213238 487798 213382
rect 487598 213210 487798 213238
rect 436200 213143 436600 213151
rect 534518 213154 534929 213538
rect 535313 213155 569529 213538
rect 569913 213155 570645 213539
rect 535313 213154 570645 213155
rect 534518 213146 570645 213154
rect 86929 212766 87129 212794
rect 86929 212622 86957 212766
rect 87101 212622 87129 212766
rect 86929 212594 87129 212622
rect 89691 212735 89891 212763
rect 89691 212591 89719 212735
rect 89863 212591 89891 212735
rect 89691 212563 89891 212591
rect 99274 212715 99474 212743
rect 99274 212571 99302 212715
rect 99446 212571 99474 212715
rect 99274 212543 99474 212571
rect 102047 212740 102247 212768
rect 102047 212596 102075 212740
rect 102219 212596 102247 212740
rect 102047 212568 102247 212596
rect 112234 212750 112434 212778
rect 112234 212606 112262 212750
rect 112406 212606 112434 212750
rect 112234 212578 112434 212606
rect 115001 212775 115201 212803
rect 115001 212631 115029 212775
rect 115173 212631 115201 212775
rect 115001 212603 115201 212631
rect 124573 212740 124773 212768
rect 124573 212596 124601 212740
rect 124745 212596 124773 212740
rect 124573 212568 124773 212596
rect 127346 212731 127546 212759
rect 127346 212587 127374 212731
rect 127518 212587 127546 212731
rect 127346 212559 127546 212587
rect 137889 212727 138089 212755
rect 137889 212583 137917 212727
rect 138061 212583 138089 212727
rect 137889 212555 138089 212583
rect 140651 212747 140851 212775
rect 140651 212603 140679 212747
rect 140823 212603 140851 212747
rect 140651 212575 140851 212603
rect 150231 212688 150431 212716
rect 150231 212544 150259 212688
rect 150403 212544 150431 212688
rect 150231 212516 150431 212544
rect 152989 212704 153189 212732
rect 152989 212560 153017 212704
rect 153161 212560 153189 212704
rect 152989 212532 153189 212560
rect 163531 212705 163731 212733
rect 163531 212561 163559 212705
rect 163703 212561 163731 212705
rect 163531 212533 163731 212561
rect 166302 212693 166502 212721
rect 166302 212549 166330 212693
rect 166474 212549 166502 212693
rect 166302 212521 166502 212549
rect 175881 212712 176081 212740
rect 175881 212568 175909 212712
rect 176053 212568 176081 212712
rect 175881 212540 176081 212568
rect 178642 212693 178842 212721
rect 178642 212549 178670 212693
rect 178814 212549 178842 212693
rect 178642 212521 178842 212549
rect 189185 212719 189385 212747
rect 189185 212575 189213 212719
rect 189357 212575 189385 212719
rect 189185 212547 189385 212575
rect 191952 212719 192152 212747
rect 191952 212575 191980 212719
rect 192124 212575 192152 212719
rect 191952 212547 192152 212575
rect 201526 212729 201726 212757
rect 214834 212749 215034 212777
rect 201526 212585 201554 212729
rect 201698 212585 201726 212729
rect 201526 212557 201726 212585
rect 204292 212707 204492 212735
rect 204292 212563 204320 212707
rect 204464 212563 204492 212707
rect 214834 212605 214862 212749
rect 215006 212605 215034 212749
rect 214834 212577 215034 212605
rect 217598 212745 217798 212773
rect 217598 212601 217626 212745
rect 217770 212601 217798 212745
rect 217598 212573 217798 212601
rect 227185 212738 227385 212766
rect 227185 212594 227213 212738
rect 227357 212594 227385 212738
rect 227185 212566 227385 212594
rect 229944 212716 230144 212744
rect 229944 212572 229972 212716
rect 230116 212572 230144 212716
rect 204292 212535 204492 212563
rect 229944 212544 230144 212572
rect 240486 212737 240686 212765
rect 240486 212593 240514 212737
rect 240658 212593 240686 212737
rect 240486 212565 240686 212593
rect 243247 212746 243447 212774
rect 332544 212770 332744 212798
rect 243247 212602 243275 212746
rect 243419 212602 243447 212746
rect 243247 212574 243447 212602
rect 252832 212727 253032 212755
rect 252832 212583 252860 212727
rect 253004 212583 253032 212727
rect 252832 212555 253032 212583
rect 255592 212727 255792 212755
rect 255592 212583 255620 212727
rect 255764 212583 255792 212727
rect 278477 212708 278677 212736
rect 268900 212677 269100 212705
rect 255592 212555 255792 212583
rect 266133 212643 266333 212671
rect 266133 212499 266161 212643
rect 266305 212499 266333 212643
rect 268900 212533 268928 212677
rect 269072 212533 269100 212677
rect 278477 212564 278505 212708
rect 278649 212564 278677 212708
rect 278477 212536 278677 212564
rect 281245 212718 281445 212746
rect 281245 212574 281273 212718
rect 281417 212574 281445 212718
rect 281245 212546 281445 212574
rect 291785 212652 291985 212680
rect 268900 212505 269100 212533
rect 291785 212508 291813 212652
rect 291957 212508 291985 212652
rect 266133 212471 266333 212499
rect 291785 212480 291985 212508
rect 294548 212673 294748 212701
rect 294548 212529 294576 212673
rect 294720 212529 294748 212673
rect 294548 212501 294748 212529
rect 304137 212693 304337 212721
rect 304137 212549 304165 212693
rect 304309 212549 304337 212693
rect 304137 212521 304337 212549
rect 306901 212688 307101 212716
rect 306901 212544 306929 212688
rect 307073 212544 307101 212688
rect 306901 212516 307101 212544
rect 317440 212708 317640 212736
rect 317440 212564 317468 212708
rect 317612 212564 317640 212708
rect 317440 212536 317640 212564
rect 320198 212708 320398 212736
rect 320198 212564 320226 212708
rect 320370 212564 320398 212708
rect 320198 212536 320398 212564
rect 329781 212735 329981 212763
rect 329781 212591 329809 212735
rect 329953 212591 329981 212735
rect 332544 212626 332572 212770
rect 332716 212626 332744 212770
rect 332544 212598 332744 212626
rect 343087 212706 343287 212734
rect 329781 212563 329981 212591
rect 343087 212562 343115 212706
rect 343259 212562 343287 212706
rect 343087 212534 343287 212562
rect 345849 212711 346049 212739
rect 345849 212567 345877 212711
rect 346021 212567 346049 212711
rect 345849 212539 346049 212567
rect 355428 212702 355628 212730
rect 355428 212558 355456 212702
rect 355600 212558 355628 212702
rect 355428 212530 355628 212558
rect 358194 212721 358394 212749
rect 358194 212577 358222 212721
rect 358366 212577 358394 212721
rect 358194 212549 358394 212577
rect 368737 212688 368937 212716
rect 368737 212544 368765 212688
rect 368909 212544 368937 212688
rect 368737 212516 368937 212544
rect 371499 212712 371699 212740
rect 371499 212568 371527 212712
rect 371671 212568 371699 212712
rect 371499 212540 371699 212568
rect 381081 212735 381281 212763
rect 381081 212591 381109 212735
rect 381253 212591 381281 212735
rect 381081 212563 381281 212591
rect 383846 212754 384046 212782
rect 383846 212610 383874 212754
rect 384018 212610 384046 212754
rect 397149 212749 397349 212777
rect 383846 212582 384046 212610
rect 394388 212699 394588 212727
rect 394388 212555 394416 212699
rect 394560 212555 394588 212699
rect 397149 212605 397177 212749
rect 397321 212605 397349 212749
rect 397149 212577 397349 212605
rect 406727 212715 406927 212743
rect 394388 212527 394588 212555
rect 406727 212571 406755 212715
rect 406899 212571 406927 212715
rect 406727 212543 406927 212571
rect 409496 212735 409696 212763
rect 409496 212591 409524 212735
rect 409668 212591 409696 212735
rect 409496 212563 409696 212591
rect 420037 212740 420237 212768
rect 420037 212596 420065 212740
rect 420209 212596 420237 212740
rect 420037 212568 420237 212596
rect 422800 212758 423000 212786
rect 422800 212614 422828 212758
rect 422972 212614 423000 212758
rect 422800 212586 423000 212614
rect 432386 212755 432586 212783
rect 432386 212611 432414 212755
rect 432558 212611 432586 212755
rect 432386 212583 432586 212611
rect 435145 212727 435345 212755
rect 435145 212583 435173 212727
rect 435317 212583 435345 212727
rect 448449 212726 448649 212754
rect 435145 212555 435345 212583
rect 445681 212672 445881 212700
rect 445681 212528 445709 212672
rect 445853 212528 445881 212672
rect 448449 212582 448477 212726
rect 448621 212582 448649 212726
rect 460793 212719 460993 212747
rect 486447 212723 486647 212751
rect 448449 212554 448649 212582
rect 458031 212687 458231 212715
rect 445681 212500 445881 212528
rect 458031 212543 458059 212687
rect 458203 212543 458231 212687
rect 460793 212575 460821 212719
rect 460965 212575 460993 212719
rect 474100 212695 474300 212723
rect 460793 212547 460993 212575
rect 471328 212641 471528 212669
rect 458031 212515 458231 212543
rect 471328 212497 471356 212641
rect 471500 212497 471528 212641
rect 474100 212551 474128 212695
rect 474272 212551 474300 212695
rect 474100 212523 474300 212551
rect 483684 212653 483884 212681
rect 471328 212469 471528 212497
rect 483684 212509 483712 212653
rect 483856 212509 483884 212653
rect 486447 212579 486475 212723
rect 486619 212579 486647 212723
rect 486447 212551 486647 212579
rect 483684 212481 483884 212509
rect -800 207380 3609 207780
rect 101200 212328 101300 212366
rect 101200 212272 101222 212328
rect 101278 212272 101300 212328
rect -800 204888 1660 207380
rect 101200 198449 101300 212272
rect 126513 212315 126613 212350
rect 126513 212259 126535 212315
rect 126591 212259 126613 212315
rect 126513 199590 126613 212259
rect 152164 212314 152264 212346
rect 152164 212258 152186 212314
rect 152242 212258 152264 212314
rect 152164 200253 152264 212258
rect 177802 212332 177902 212346
rect 177802 212310 177903 212332
rect 177802 212254 177825 212310
rect 177881 212254 177903 212310
rect 177802 212232 177903 212254
rect 203459 212316 203559 212347
rect 229099 212338 229199 212350
rect 203459 212260 203481 212316
rect 203537 212260 203559 212316
rect 177802 201219 177902 212232
rect 203459 202152 203559 212260
rect 229098 212316 229199 212338
rect 229098 212260 229120 212316
rect 229176 212260 229199 212316
rect 229098 212238 229199 212260
rect 229099 202919 229199 212238
rect 254765 212313 254865 212346
rect 254765 212257 254787 212313
rect 254843 212257 254865 212313
rect 254765 203441 254865 212257
rect 280408 212316 280508 212346
rect 306062 212333 306162 212347
rect 280408 212260 280430 212316
rect 280486 212260 280508 212316
rect 280408 204373 280508 212260
rect 306061 212311 306162 212333
rect 306061 212255 306083 212311
rect 306139 212255 306162 212311
rect 306061 212233 306162 212255
rect 306062 205676 306162 212233
rect 331707 212311 331807 212342
rect 331707 212255 331729 212311
rect 331785 212255 331807 212311
rect 331707 206532 331807 212255
rect 357354 212320 357454 212346
rect 357354 212264 357376 212320
rect 357432 212264 357454 212320
rect 357354 207292 357454 212264
rect 382989 212316 383089 212342
rect 382989 212260 383011 212316
rect 383067 212260 383089 212316
rect 382989 207949 383089 212260
rect 408655 212316 408755 212348
rect 408655 212260 408677 212316
rect 408733 212260 408755 212316
rect 408655 209166 408755 212260
rect 434292 212311 434392 212344
rect 434292 212255 434314 212311
rect 434370 212255 434392 212311
rect 434292 209736 434392 212255
rect 459957 212312 460057 212341
rect 459957 212256 459979 212312
rect 460035 212256 460057 212312
rect 459957 210252 460057 212256
rect 485597 212336 485697 212347
rect 485597 212314 485698 212336
rect 485597 212258 485620 212314
rect 485676 212258 485698 212314
rect 485597 212236 485698 212258
rect 485597 210971 485697 212236
rect 485597 210871 537813 210971
rect 459957 210152 537114 210252
rect 434292 209636 536608 209736
rect 408655 209066 535695 209166
rect 382989 207849 534858 207949
rect 357354 207192 534392 207292
rect 331707 206432 533822 206532
rect 306062 205576 533014 205676
rect 280408 204273 532182 204373
rect 254765 203341 531647 203441
rect 229099 202819 531015 202919
rect 203459 202052 530388 202152
rect 177802 201119 529418 201219
rect 152164 200153 528694 200253
rect 126513 199490 528117 199590
rect 101200 198349 527487 198449
rect 484635 197100 526534 197122
rect 484635 197044 484658 197100
rect 484714 197044 526534 197100
rect 484635 197022 526534 197044
rect 458986 195926 525631 195948
rect 458986 195870 459011 195926
rect 459067 195870 525631 195926
rect 458986 195848 525631 195870
rect 433348 194511 523042 194533
rect 433348 194455 433370 194511
rect 433426 194455 523042 194511
rect 433348 194433 523042 194455
rect 407692 192377 521310 192399
rect 407692 192321 407725 192377
rect 407781 192321 521310 192377
rect 407692 192299 521310 192321
rect 100236 192094 100336 192116
rect 100236 192038 100258 192094
rect 100314 192038 100336 192094
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 241 124905 441 124937
rect 241 124888 273 124905
rect -800 124776 273 124888
rect 241 124769 273 124776
rect 409 124888 441 124905
rect 409 124776 480 124888
rect 409 124769 441 124776
rect 241 124737 441 124769
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 100236 92874 100336 192038
rect 125541 191931 125641 191953
rect 125541 191930 125563 191931
rect 125540 191875 125563 191930
rect 125619 191875 125641 191931
rect 125540 191853 125641 191875
rect 125540 140377 125640 191853
rect 382031 191030 520181 191052
rect 382031 190974 382053 191030
rect 382109 190974 520181 191030
rect 382031 190952 520181 190974
rect 176840 190325 176940 190380
rect 176840 190269 176862 190325
rect 176918 190269 176940 190325
rect 102885 140277 125640 140377
rect 151197 189955 151297 189977
rect 151197 189899 151219 189955
rect 151275 189899 151297 189955
rect 102885 95212 102985 140277
rect 151197 136071 151297 189899
rect 106298 135971 151297 136071
rect 106298 97995 106398 135971
rect 176840 132329 176940 190269
rect 356393 189652 519194 189674
rect 356393 189596 356415 189652
rect 356471 189596 519194 189652
rect 356393 189574 519194 189596
rect 253784 188715 253884 188737
rect 253784 188659 253806 188715
rect 253862 188659 253884 188715
rect 253784 188637 253884 188659
rect 108268 132229 176940 132329
rect 202478 188135 202578 188140
rect 202478 188113 202579 188135
rect 202478 188057 202501 188113
rect 202557 188057 202579 188113
rect 202478 188035 202579 188057
rect 108268 99423 108368 132229
rect 202478 129958 202578 188035
rect 110027 129858 202578 129958
rect 228146 187406 228246 187447
rect 228146 187350 228168 187406
rect 228224 187350 228246 187406
rect 110027 100560 110127 129858
rect 228146 126832 228246 187350
rect 111540 126732 228246 126832
rect 111540 101575 111640 126732
rect 253784 123611 253884 187468
rect 330739 187409 517284 187431
rect 330739 187353 330761 187409
rect 330817 187353 517284 187409
rect 330739 187331 517284 187353
rect 113906 123511 253884 123611
rect 279438 186937 279538 187000
rect 279438 186881 279460 186937
rect 279516 186881 279538 186937
rect 113906 102702 114006 123511
rect 279438 120513 279538 186881
rect 305089 186372 515989 186394
rect 305089 186316 305111 186372
rect 305167 186316 515989 186372
rect 305089 186294 515989 186316
rect 114934 120413 279538 120513
rect 114934 104098 115034 120413
rect 114934 103998 377791 104098
rect 377585 103392 377685 103414
rect 377585 103336 377607 103392
rect 377663 103336 377685 103392
rect 377585 103314 377685 103336
rect 113906 102680 375143 102702
rect 113906 102624 374062 102680
rect 374118 102624 375143 102680
rect 113906 102602 375143 102624
rect 111540 101553 370678 101575
rect 111540 101497 370515 101553
rect 370571 101497 370678 101553
rect 111540 101475 370678 101497
rect 110027 100538 367137 100560
rect 110027 100482 366968 100538
rect 367024 100482 367137 100538
rect 110027 100460 367137 100482
rect 108268 99401 363579 99423
rect 108268 99345 363423 99401
rect 363479 99345 363579 99401
rect 108268 99323 363579 99345
rect 359855 97995 359955 97996
rect 106298 97974 360063 97995
rect 106298 97918 359877 97974
rect 359933 97918 360063 97974
rect 106298 97895 360063 97918
rect 356322 95212 356422 95213
rect 102885 95191 356513 95212
rect 102885 95135 356344 95191
rect 356400 95135 356513 95191
rect 102885 95112 356513 95135
rect 100236 92852 352941 92874
rect 100236 92796 352774 92852
rect 352830 92796 352941 92852
rect 100236 92774 352941 92796
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 515889 60405 515989 186294
rect 381029 60383 515989 60405
rect 381029 60327 381143 60383
rect 381199 60327 515989 60383
rect 381029 60305 515989 60327
rect 517184 59318 517284 187331
rect 384600 59218 517284 59318
rect 519094 58452 519194 189574
rect 388163 58430 519194 58452
rect 388163 58374 388239 58430
rect 388295 58374 519194 58430
rect 388163 58352 519194 58374
rect 520081 58049 520181 190952
rect 391626 58027 520181 58049
rect 391626 57971 391787 58027
rect 391843 57971 520181 58027
rect 391626 57949 520181 57971
rect 521210 57722 521310 192299
rect 395265 57700 521310 57722
rect 395265 57644 395335 57700
rect 395391 57644 521310 57700
rect 395265 57622 521310 57644
rect 522942 57072 523042 194433
rect 398743 57050 523042 57072
rect 398743 56994 398880 57050
rect 398936 56994 523042 57050
rect 398743 56972 523042 56994
rect 525531 56570 525631 195848
rect 402266 56548 525631 56570
rect 402266 56492 402422 56548
rect 402478 56492 525631 56548
rect 402266 56470 525631 56492
rect 526434 56055 526534 197022
rect 405879 56033 526534 56055
rect 405879 55977 405983 56033
rect 406039 55977 526534 56033
rect 405879 55955 526534 55977
rect 527387 54187 527487 198349
rect 409408 54165 527487 54187
rect 409408 54109 409531 54165
rect 409587 54109 527487 54165
rect 409408 54087 527487 54109
rect 528017 53371 528117 199490
rect 412965 53349 528117 53371
rect 412965 53293 413076 53349
rect 413132 53293 528117 53349
rect 412965 53271 528117 53293
rect 528594 52794 528694 200153
rect 416521 52772 528694 52794
rect 416521 52716 416628 52772
rect 416684 52716 528694 52772
rect 416521 52694 528694 52716
rect 529318 52272 529418 201119
rect 420063 52250 529418 52272
rect 420063 52194 420154 52250
rect 420210 52194 529418 52250
rect 420063 52172 529418 52194
rect 530288 51935 530388 202052
rect 423590 51913 530388 51935
rect 423590 51857 423714 51913
rect 423770 51857 530388 51913
rect 423590 51835 530388 51857
rect 530915 50936 531015 202819
rect 427146 50914 531015 50936
rect 427146 50858 427266 50914
rect 427322 50858 531015 50914
rect 427146 50836 531015 50858
rect 531547 50379 531647 203341
rect 430679 50357 531647 50379
rect 430679 50301 430790 50357
rect 430846 50301 531647 50357
rect 430679 50279 531647 50301
rect 532082 49436 532182 204273
rect 434213 49414 532182 49436
rect 434213 49358 434349 49414
rect 434405 49358 532182 49414
rect 434213 49336 532182 49358
rect 532914 48782 533014 205576
rect 437774 48760 533014 48782
rect 437774 48704 437875 48760
rect 437931 48704 533014 48760
rect 437774 48682 533014 48704
rect 533722 48117 533822 206432
rect 441239 48095 533822 48117
rect 441239 48039 441438 48095
rect 441494 48039 533822 48095
rect 441239 48017 533822 48039
rect 534292 47475 534392 207192
rect 444904 47453 534392 47475
rect 444904 47397 444991 47453
rect 445047 47397 534392 47453
rect 444904 47375 534392 47397
rect 534758 46947 534858 207849
rect 448393 46925 534858 46947
rect 448393 46869 448515 46925
rect 448571 46869 534858 46925
rect 448393 46847 534858 46869
rect 535595 46583 535695 209066
rect 451958 46561 535695 46583
rect 451958 46505 452075 46561
rect 452131 46505 535695 46561
rect 451958 46483 535695 46505
rect 536508 45736 536608 209636
rect 455519 45714 536608 45736
rect 455519 45658 455623 45714
rect 455679 45658 536608 45714
rect 455519 45636 536608 45658
rect 537014 45179 537114 210152
rect 459048 45157 537114 45179
rect 459048 45101 459169 45157
rect 459225 45101 537114 45157
rect 459048 45079 537114 45101
rect 537713 44484 537813 210871
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 582340 149156 584800 151630
rect 578061 148956 584800 149156
rect 578061 145751 578261 148956
rect 582340 146830 584800 148956
rect 568794 144895 578985 145751
rect 568794 144511 570135 144895
rect 570519 144511 578985 144895
rect 568794 143351 578985 144511
rect 577901 139226 578301 143351
rect 582340 139226 584800 141630
rect 577901 138826 584800 139226
rect 582340 136830 584800 138826
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 462616 44462 537813 44484
rect 462616 44406 462719 44462
rect 462775 44406 537813 44462
rect 462616 44384 537813 44406
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 583220 500050 583318 500162
rect 660 462398 780 462510
rect 583180 455628 583296 455740
rect 676 419176 738 419288
<< via3 >>
rect 95445 687797 95829 687801
rect 95445 687421 95449 687797
rect 95449 687421 95825 687797
rect 95825 687421 95829 687797
rect 95445 687417 95829 687421
rect 120770 687611 121154 687615
rect 120770 687235 120774 687611
rect 120774 687235 121150 687611
rect 121150 687235 121154 687611
rect 120770 687231 121154 687235
rect 146427 687489 146811 687493
rect 146427 687113 146431 687489
rect 146431 687113 146807 687489
rect 146807 687113 146811 687489
rect 146427 687109 146811 687113
rect 172228 688020 172612 688024
rect 172228 687644 172232 688020
rect 172232 687644 172608 688020
rect 172608 687644 172612 688020
rect 172228 687640 172612 687644
rect 216366 687580 216750 687584
rect 216366 687204 216370 687580
rect 216370 687204 216746 687580
rect 216746 687204 216750 687580
rect 216366 687200 216750 687204
rect 223347 687655 223731 687659
rect 223347 687279 223351 687655
rect 223351 687279 223727 687655
rect 223727 687279 223731 687655
rect 223347 687275 223731 687279
rect 249017 687558 249401 687562
rect 249017 687182 249021 687558
rect 249021 687182 249397 687558
rect 249397 687182 249401 687558
rect 249017 687178 249401 687182
rect 274686 687574 275070 687578
rect 274686 687198 274690 687574
rect 274690 687198 275066 687574
rect 275066 687198 275070 687574
rect 274686 687194 275070 687198
rect 300311 687610 300695 687614
rect 300311 687234 300315 687610
rect 300315 687234 300691 687610
rect 300691 687234 300695 687610
rect 300311 687230 300695 687234
rect 325947 687575 326331 687579
rect 325947 687199 325951 687575
rect 325951 687199 326327 687575
rect 326327 687199 326331 687575
rect 325947 687195 326331 687199
rect 351612 687557 351996 687561
rect 351612 687181 351616 687557
rect 351616 687181 351992 687557
rect 351992 687181 351996 687557
rect 351612 687177 351996 687181
rect 377273 687519 377657 687523
rect 377273 687143 377277 687519
rect 377277 687143 377653 687519
rect 377653 687143 377657 687519
rect 377273 687139 377657 687143
rect 412449 687636 412833 687640
rect 412449 687260 412453 687636
rect 412453 687260 412829 687636
rect 412829 687260 412833 687636
rect 412449 687256 412833 687260
rect 428575 687626 428959 687630
rect 428575 687250 428579 687626
rect 428579 687250 428955 687626
rect 428955 687250 428959 687626
rect 428575 687246 428959 687250
rect 454209 687695 454593 687699
rect 454209 687319 454213 687695
rect 454213 687319 454589 687695
rect 454589 687319 454593 687695
rect 454209 687315 454593 687319
rect 479858 687701 480242 687705
rect 479858 687325 479862 687701
rect 479862 687325 480238 687701
rect 480238 687325 480242 687701
rect 479858 687321 480242 687325
rect 512525 687670 513309 688454
rect 522690 687712 523474 688496
rect 560582 639792 566726 644576
rect 560582 629792 566726 634576
rect 556255 550570 562319 555354
rect 37859 542707 38243 542711
rect 37859 542331 37863 542707
rect 37863 542331 38239 542707
rect 38239 542331 38243 542707
rect 37859 542327 38243 542331
rect 556255 540570 562319 545354
rect 10434 530632 10818 531016
rect 569788 530633 570172 531017
rect 76152 438023 76296 438027
rect 76152 437887 76156 438023
rect 76156 437887 76292 438023
rect 76292 437887 76296 438023
rect 76152 437883 76296 437887
rect 76169 435267 76313 435271
rect 76169 435131 76173 435267
rect 76173 435131 76309 435267
rect 76309 435131 76313 435267
rect 76169 435127 76313 435131
rect 77100 434111 77244 434115
rect 77100 433975 77104 434111
rect 77104 433975 77240 434111
rect 77240 433975 77244 434111
rect 77100 433971 77244 433975
rect 79031 433163 79175 433167
rect 79031 433027 79035 433163
rect 79035 433027 79171 433163
rect 79171 433027 79175 433163
rect 79031 433023 79175 433027
rect 76179 424683 76323 424687
rect 76179 424547 76183 424683
rect 76183 424547 76319 424683
rect 76319 424547 76323 424683
rect 76179 424543 76323 424547
rect 76194 421917 76338 421921
rect 76194 421781 76198 421917
rect 76198 421781 76334 421917
rect 76334 421781 76338 421917
rect 76194 421777 76338 421781
rect 77133 420759 77277 420763
rect 77133 420623 77137 420759
rect 77137 420623 77273 420759
rect 77273 420623 77277 420759
rect 77133 420619 77277 420623
rect 79022 419816 79166 419820
rect 79022 419680 79026 419816
rect 79026 419680 79162 419816
rect 79162 419680 79166 419816
rect 79022 419676 79166 419680
rect 76163 411339 76307 411343
rect 76163 411203 76167 411339
rect 76167 411203 76303 411339
rect 76303 411203 76307 411339
rect 76163 411199 76307 411203
rect 76194 408572 76338 408576
rect 76194 408436 76198 408572
rect 76198 408436 76334 408572
rect 76334 408436 76338 408572
rect 76194 408432 76338 408436
rect 77121 407419 77265 407423
rect 77121 407283 77125 407419
rect 77125 407283 77261 407419
rect 77261 407283 77265 407419
rect 77121 407279 77265 407283
rect 79006 406471 79150 406475
rect 79006 406335 79010 406471
rect 79010 406335 79146 406471
rect 79146 406335 79150 406471
rect 79006 406331 79150 406335
rect 76176 397984 76320 397988
rect 76176 397848 76180 397984
rect 76180 397848 76316 397984
rect 76316 397848 76320 397984
rect 76176 397844 76320 397848
rect 76181 395230 76325 395234
rect 76181 395094 76185 395230
rect 76185 395094 76321 395230
rect 76321 395094 76325 395230
rect 76181 395090 76325 395094
rect 77133 394070 77277 394074
rect 77133 393934 77137 394070
rect 77137 393934 77273 394070
rect 77273 393934 77277 394070
rect 77133 393930 77277 393934
rect 79031 393131 79175 393135
rect 79031 392995 79035 393131
rect 79035 392995 79171 393131
rect 79171 392995 79175 393131
rect 79031 392991 79175 392995
rect 76151 384644 76295 384648
rect 76151 384508 76155 384644
rect 76155 384508 76291 384644
rect 76291 384508 76295 384644
rect 76151 384504 76295 384508
rect 76156 381882 76300 381886
rect 76156 381746 76160 381882
rect 76160 381746 76296 381882
rect 76296 381746 76300 381882
rect 76156 381742 76300 381746
rect 77121 380726 77265 380730
rect 77121 380590 77125 380726
rect 77125 380590 77261 380726
rect 77261 380590 77265 380726
rect 77121 380586 77265 380590
rect 78997 379784 79141 379788
rect 78997 379648 79001 379784
rect 79001 379648 79137 379784
rect 79137 379648 79141 379784
rect 78997 379644 79141 379648
rect 76171 371302 76315 371306
rect 76171 371166 76175 371302
rect 76175 371166 76311 371302
rect 76311 371166 76315 371302
rect 76171 371162 76315 371166
rect 76174 368541 76318 368545
rect 76174 368405 76178 368541
rect 76178 368405 76314 368541
rect 76314 368405 76318 368541
rect 76174 368401 76318 368405
rect 77083 367381 77227 367385
rect 77083 367245 77087 367381
rect 77087 367245 77223 367381
rect 77223 367245 77227 367381
rect 77083 367241 77227 367245
rect 79016 366435 79160 366439
rect 79016 366299 79020 366435
rect 79020 366299 79156 366435
rect 79156 366299 79160 366435
rect 79016 366295 79160 366299
rect 76161 357953 76305 357957
rect 76161 357817 76165 357953
rect 76165 357817 76301 357953
rect 76301 357817 76305 357953
rect 76161 357813 76305 357817
rect 76181 355196 76325 355200
rect 76181 355060 76185 355196
rect 76185 355060 76321 355196
rect 76321 355060 76325 355196
rect 76181 355056 76325 355060
rect 77173 354037 77317 354041
rect 77173 353901 77177 354037
rect 77177 353901 77313 354037
rect 77313 353901 77317 354037
rect 77173 353897 77317 353901
rect 79020 353095 79164 353099
rect 79020 352959 79024 353095
rect 79024 352959 79160 353095
rect 79160 352959 79164 353095
rect 79020 352955 79164 352959
rect 76128 344608 76272 344612
rect 76128 344472 76132 344608
rect 76132 344472 76268 344608
rect 76268 344472 76272 344608
rect 76128 344468 76272 344472
rect 76151 341846 76295 341850
rect 76151 341710 76155 341846
rect 76155 341710 76291 341846
rect 76291 341710 76295 341846
rect 76151 341706 76295 341710
rect 77139 340695 77283 340699
rect 77139 340559 77143 340695
rect 77143 340559 77279 340695
rect 77279 340559 77283 340695
rect 77139 340555 77283 340559
rect 79027 339746 79171 339750
rect 79027 339610 79031 339746
rect 79031 339610 79167 339746
rect 79167 339610 79171 339746
rect 79027 339606 79171 339610
rect 76171 331264 76315 331268
rect 76171 331128 76175 331264
rect 76175 331128 76311 331264
rect 76311 331128 76315 331264
rect 76171 331124 76315 331128
rect 76175 328506 76319 328510
rect 76175 328370 76179 328506
rect 76179 328370 76315 328506
rect 76315 328370 76319 328506
rect 76175 328366 76319 328370
rect 77127 327352 77271 327356
rect 77127 327216 77131 327352
rect 77131 327216 77267 327352
rect 77267 327216 77271 327352
rect 77127 327212 77271 327216
rect 79039 326398 79183 326402
rect 79039 326262 79043 326398
rect 79043 326262 79179 326398
rect 79179 326262 79183 326398
rect 79039 326258 79183 326262
rect 76183 317912 76327 317916
rect 76183 317776 76187 317912
rect 76187 317776 76323 317912
rect 76323 317776 76327 317912
rect 76183 317772 76327 317776
rect 76171 315161 76315 315165
rect 76171 315025 76175 315161
rect 76175 315025 76311 315161
rect 76311 315025 76315 315161
rect 76171 315021 76315 315025
rect 77132 314006 77276 314010
rect 77132 313870 77136 314006
rect 77136 313870 77272 314006
rect 77272 313870 77276 314006
rect 77132 313866 77276 313870
rect 78998 313060 79142 313064
rect 78998 312924 79002 313060
rect 79002 312924 79138 313060
rect 79138 312924 79142 313060
rect 78998 312920 79142 312924
rect 76166 304571 76310 304575
rect 76166 304435 76170 304571
rect 76170 304435 76306 304571
rect 76306 304435 76310 304571
rect 76166 304431 76310 304435
rect 76181 301814 76325 301818
rect 76181 301678 76185 301814
rect 76185 301678 76321 301814
rect 76321 301678 76325 301814
rect 76181 301674 76325 301678
rect 77138 300655 77282 300659
rect 77138 300519 77142 300655
rect 77142 300519 77278 300655
rect 77278 300519 77282 300655
rect 77138 300515 77282 300519
rect 79011 299709 79155 299713
rect 79011 299573 79015 299709
rect 79015 299573 79151 299709
rect 79151 299573 79155 299709
rect 79011 299569 79155 299573
rect 76166 291231 76310 291235
rect 76166 291095 76170 291231
rect 76170 291095 76306 291231
rect 76306 291095 76310 291231
rect 76166 291091 76310 291095
rect 76156 288478 76300 288482
rect 76156 288342 76160 288478
rect 76160 288342 76296 288478
rect 76296 288342 76300 288478
rect 76156 288338 76300 288342
rect 77135 287312 77279 287316
rect 77135 287176 77139 287312
rect 77139 287176 77275 287312
rect 77275 287176 77279 287312
rect 77135 287172 77279 287176
rect 79009 286366 79153 286370
rect 79009 286230 79013 286366
rect 79013 286230 79149 286366
rect 79149 286230 79153 286366
rect 79009 286226 79153 286230
rect 76174 277897 76318 277901
rect 76174 277761 76178 277897
rect 76178 277761 76314 277897
rect 76314 277761 76318 277897
rect 76174 277757 76318 277761
rect 76174 275119 76318 275123
rect 76174 274983 76178 275119
rect 76178 274983 76314 275119
rect 76314 274983 76318 275119
rect 76174 274979 76318 274983
rect 77146 273968 77290 273972
rect 77146 273832 77150 273968
rect 77150 273832 77286 273968
rect 77286 273832 77290 273968
rect 77146 273828 77290 273832
rect 79016 273027 79160 273031
rect 79016 272891 79020 273027
rect 79020 272891 79156 273027
rect 79156 272891 79160 273027
rect 79016 272887 79160 272891
rect 76185 264540 76329 264544
rect 76185 264404 76189 264540
rect 76189 264404 76325 264540
rect 76325 264404 76329 264540
rect 76185 264400 76329 264404
rect 76197 261781 76341 261785
rect 76197 261645 76201 261781
rect 76201 261645 76337 261781
rect 76337 261645 76341 261781
rect 76197 261641 76341 261645
rect 77148 260623 77292 260627
rect 77148 260487 77152 260623
rect 77152 260487 77288 260623
rect 77288 260487 77292 260623
rect 77148 260483 77292 260487
rect 79003 259676 79147 259680
rect 79003 259540 79007 259676
rect 79007 259540 79143 259676
rect 79143 259540 79147 259676
rect 79003 259536 79147 259540
rect 76182 251191 76326 251195
rect 76182 251055 76186 251191
rect 76186 251055 76322 251191
rect 76322 251055 76326 251191
rect 76182 251051 76326 251055
rect 76180 248432 76324 248436
rect 76180 248296 76184 248432
rect 76184 248296 76320 248432
rect 76320 248296 76324 248432
rect 76180 248292 76324 248296
rect 77126 247276 77270 247280
rect 77126 247140 77130 247276
rect 77130 247140 77266 247276
rect 77266 247140 77270 247276
rect 77126 247136 77270 247140
rect 79017 246330 79161 246334
rect 79017 246194 79021 246330
rect 79021 246194 79157 246330
rect 79157 246194 79161 246330
rect 79017 246190 79161 246194
rect 76229 237818 76373 237822
rect 76229 237682 76233 237818
rect 76233 237682 76369 237818
rect 76369 237682 76373 237818
rect 76229 237678 76373 237682
rect 76227 235050 76371 235054
rect 76227 234914 76231 235050
rect 76231 234914 76367 235050
rect 76367 234914 76371 235050
rect 76227 234910 76371 234914
rect 77104 233894 77248 233898
rect 77104 233758 77108 233894
rect 77108 233758 77244 233894
rect 77244 233758 77248 233894
rect 77104 233754 77248 233758
rect 79012 232948 79156 232952
rect 79012 232812 79016 232948
rect 79016 232812 79152 232948
rect 79152 232812 79156 232948
rect 79012 232808 79156 232812
rect 539194 231700 540778 233284
rect 91818 215228 91962 215232
rect 91818 215092 91822 215228
rect 91822 215092 91958 215228
rect 91958 215092 91962 215228
rect 91818 215088 91962 215092
rect 104163 215219 104307 215223
rect 104163 215083 104167 215219
rect 104167 215083 104303 215219
rect 104303 215083 104307 215219
rect 104163 215079 104307 215083
rect 117137 215241 117281 215245
rect 117137 215105 117141 215241
rect 117141 215105 117277 215241
rect 117277 215105 117281 215241
rect 117137 215101 117281 215105
rect 129472 215179 129616 215183
rect 129472 215043 129476 215179
rect 129476 215043 129612 215179
rect 129612 215043 129616 215179
rect 129472 215039 129616 215043
rect 142787 215195 142931 215199
rect 142787 215059 142791 215195
rect 142791 215059 142927 215195
rect 142927 215059 142931 215195
rect 142787 215055 142931 215059
rect 155127 215225 155271 215229
rect 155127 215089 155131 215225
rect 155131 215089 155267 215225
rect 155267 215089 155271 215225
rect 155127 215085 155271 215089
rect 168429 215182 168573 215186
rect 168429 215046 168433 215182
rect 168433 215046 168569 215182
rect 168569 215046 168573 215182
rect 168429 215042 168573 215046
rect 180783 215213 180927 215217
rect 180783 215077 180787 215213
rect 180787 215077 180923 215213
rect 180923 215077 180927 215213
rect 180783 215073 180927 215077
rect 194072 215241 194216 215245
rect 194072 215105 194076 215241
rect 194076 215105 194212 215241
rect 194212 215105 194216 215241
rect 194072 215101 194216 215105
rect 206430 215219 206574 215223
rect 206430 215083 206434 215219
rect 206434 215083 206570 215219
rect 206570 215083 206574 215219
rect 206430 215079 206574 215083
rect 219727 215218 219871 215222
rect 219727 215082 219731 215218
rect 219731 215082 219867 215218
rect 219867 215082 219871 215218
rect 219727 215078 219871 215082
rect 232074 215253 232218 215257
rect 232074 215117 232078 215253
rect 232078 215117 232214 215253
rect 232214 215117 232218 215253
rect 232074 215113 232218 215117
rect 245378 215237 245522 215241
rect 245378 215101 245382 215237
rect 245382 215101 245518 215237
rect 245518 215101 245522 215237
rect 245378 215097 245522 215101
rect 257723 215268 257867 215272
rect 257723 215132 257727 215268
rect 257727 215132 257863 215268
rect 257863 215132 257867 215268
rect 257723 215128 257867 215132
rect 271032 215249 271176 215253
rect 271032 215113 271036 215249
rect 271036 215113 271172 215249
rect 271172 215113 271176 215249
rect 271032 215109 271176 215113
rect 283375 215231 283519 215235
rect 283375 215095 283379 215231
rect 283379 215095 283515 215231
rect 283515 215095 283519 215231
rect 283375 215091 283519 215095
rect 296678 215227 296822 215231
rect 296678 215091 296682 215227
rect 296682 215091 296818 215227
rect 296818 215091 296822 215227
rect 296678 215087 296822 215091
rect 309022 215234 309166 215238
rect 309022 215098 309026 215234
rect 309026 215098 309162 215234
rect 309162 215098 309166 215234
rect 309022 215094 309166 215098
rect 322329 215211 322473 215215
rect 322329 215075 322333 215211
rect 322333 215075 322469 215211
rect 322469 215075 322473 215211
rect 322329 215071 322473 215075
rect 334673 215241 334817 215245
rect 334673 215105 334677 215241
rect 334677 215105 334813 215241
rect 334813 215105 334817 215241
rect 334673 215101 334817 215105
rect 347979 215211 348123 215215
rect 347979 215075 347983 215211
rect 347983 215075 348119 215211
rect 348119 215075 348123 215211
rect 347979 215071 348123 215075
rect 360323 215223 360467 215227
rect 360323 215087 360327 215223
rect 360327 215087 360463 215223
rect 360463 215087 360467 215223
rect 360323 215083 360467 215087
rect 373628 215215 373772 215219
rect 373628 215079 373632 215215
rect 373632 215079 373768 215215
rect 373768 215079 373772 215215
rect 373628 215075 373772 215079
rect 385973 215242 386117 215246
rect 385973 215106 385977 215242
rect 385977 215106 386113 215242
rect 386113 215106 386117 215242
rect 385973 215102 386117 215106
rect 399278 215241 399422 215245
rect 399278 215105 399282 215241
rect 399282 215105 399418 215241
rect 399418 215105 399422 215241
rect 399278 215101 399422 215105
rect 411627 215207 411771 215211
rect 411627 215071 411631 215207
rect 411631 215071 411767 215207
rect 411767 215071 411771 215207
rect 411627 215067 411771 215071
rect 424927 215210 425071 215214
rect 424927 215074 424931 215210
rect 424931 215074 425067 215210
rect 425067 215074 425071 215210
rect 424927 215070 425071 215074
rect 437275 215228 437419 215232
rect 437275 215092 437279 215228
rect 437279 215092 437415 215228
rect 437415 215092 437419 215228
rect 437275 215088 437419 215092
rect 450571 215228 450715 215232
rect 450571 215092 450575 215228
rect 450575 215092 450711 215228
rect 450711 215092 450715 215228
rect 450571 215088 450715 215092
rect 462922 215215 463066 215219
rect 462922 215079 462926 215215
rect 462926 215079 463062 215215
rect 463062 215079 463066 215215
rect 462922 215075 463066 215079
rect 476234 215203 476378 215207
rect 476234 215067 476238 215203
rect 476238 215067 476374 215203
rect 476374 215067 476378 215203
rect 476234 215063 476378 215067
rect 488575 215221 488719 215225
rect 488575 215085 488579 215221
rect 488579 215085 488715 215221
rect 488715 215085 488719 215221
rect 488575 215081 488719 215085
rect 9842 214527 10226 214911
rect 90871 213423 91015 213427
rect 90871 213287 90875 213423
rect 90875 213287 91011 213423
rect 91011 213287 91015 213423
rect 90871 213283 91015 213287
rect 103221 213421 103365 213425
rect 103221 213285 103225 213421
rect 103225 213285 103361 213421
rect 103361 213285 103365 213421
rect 103221 213281 103365 213285
rect 116181 213422 116325 213426
rect 116181 213286 116185 213422
rect 116185 213286 116321 213422
rect 116321 213286 116325 213422
rect 116181 213282 116325 213286
rect 128524 213381 128668 213385
rect 128524 213245 128528 213381
rect 128528 213245 128664 213381
rect 128664 213245 128668 213381
rect 128524 213241 128668 213245
rect 141829 213341 141973 213345
rect 141829 213205 141833 213341
rect 141833 213205 141969 213341
rect 141969 213205 141973 213341
rect 141829 213201 141973 213205
rect 154173 213406 154317 213410
rect 154173 213270 154177 213406
rect 154177 213270 154313 213406
rect 154313 213270 154317 213406
rect 154173 213266 154317 213270
rect 167484 213367 167628 213371
rect 167484 213231 167488 213367
rect 167488 213231 167624 213367
rect 167624 213231 167628 213367
rect 167484 213227 167628 213231
rect 179828 213401 179972 213405
rect 179828 213265 179832 213401
rect 179832 213265 179968 213401
rect 179968 213265 179972 213401
rect 179828 213261 179972 213265
rect 193138 213393 193282 213397
rect 193138 213257 193142 213393
rect 193142 213257 193278 213393
rect 193278 213257 193282 213393
rect 193138 213253 193282 213257
rect 205474 213407 205618 213411
rect 205474 213271 205478 213407
rect 205478 213271 205614 213407
rect 205614 213271 205618 213407
rect 205474 213267 205618 213271
rect 218779 213408 218923 213412
rect 218779 213272 218783 213408
rect 218783 213272 218919 213408
rect 218919 213272 218923 213408
rect 218779 213268 218923 213272
rect 231129 213395 231273 213399
rect 231129 213259 231133 213395
rect 231133 213259 231269 213395
rect 231269 213259 231273 213395
rect 231129 213255 231273 213259
rect 244428 213385 244572 213389
rect 244428 213249 244432 213385
rect 244432 213249 244568 213385
rect 244568 213249 244572 213385
rect 244428 213245 244572 213249
rect 256777 213405 256921 213409
rect 256777 213269 256781 213405
rect 256781 213269 256917 213405
rect 256917 213269 256921 213405
rect 256777 213265 256921 213269
rect 270086 213386 270230 213390
rect 270086 213250 270090 213386
rect 270090 213250 270226 213386
rect 270226 213250 270230 213386
rect 270086 213246 270230 213250
rect 282430 213363 282574 213367
rect 282430 213227 282434 213363
rect 282434 213227 282570 213363
rect 282570 213227 282574 213363
rect 282430 213223 282574 213227
rect 295733 213378 295877 213382
rect 295733 213242 295737 213378
rect 295737 213242 295873 213378
rect 295873 213242 295877 213378
rect 295733 213238 295877 213242
rect 308081 213336 308225 213340
rect 308081 213200 308085 213336
rect 308085 213200 308221 213336
rect 308221 213200 308225 213336
rect 308081 213196 308225 213200
rect 321379 213395 321523 213399
rect 321379 213259 321383 213395
rect 321383 213259 321519 213395
rect 321519 213259 321523 213395
rect 321379 213255 321523 213259
rect 333724 213352 333868 213356
rect 333724 213216 333728 213352
rect 333728 213216 333864 213352
rect 333864 213216 333868 213352
rect 333724 213212 333868 213216
rect 347030 213419 347174 213423
rect 347030 213283 347034 213419
rect 347034 213283 347170 213419
rect 347170 213283 347174 213419
rect 347030 213279 347174 213283
rect 359379 213407 359523 213411
rect 359379 213271 359383 213407
rect 359383 213271 359519 213407
rect 359519 213271 359523 213407
rect 359379 213267 359523 213271
rect 372682 213419 372826 213423
rect 372682 213283 372686 213419
rect 372686 213283 372822 213419
rect 372822 213283 372826 213419
rect 372682 213279 372826 213283
rect 385029 213420 385173 213424
rect 385029 213284 385033 213420
rect 385033 213284 385169 213420
rect 385169 213284 385173 213420
rect 385029 213280 385173 213284
rect 398326 213415 398470 213419
rect 398326 213279 398330 213415
rect 398330 213279 398466 213415
rect 398466 213279 398470 213415
rect 398326 213275 398470 213279
rect 410674 213415 410818 213419
rect 410674 213279 410678 213415
rect 410678 213279 410814 213415
rect 410814 213279 410818 213415
rect 410674 213275 410818 213279
rect 423983 213418 424127 213422
rect 423983 213282 423987 213418
rect 423987 213282 424123 213418
rect 424123 213282 424127 213418
rect 423983 213278 424127 213282
rect 436208 213531 436592 213535
rect 436208 213155 436212 213531
rect 436212 213155 436588 213531
rect 436588 213155 436592 213531
rect 436208 213151 436592 213155
rect 449633 213411 449777 213415
rect 449633 213275 449637 213411
rect 449637 213275 449773 213411
rect 449773 213275 449777 213411
rect 449633 213271 449777 213275
rect 461981 213409 462125 213413
rect 461981 213273 461985 213409
rect 461985 213273 462121 213409
rect 462121 213273 462125 213409
rect 461981 213269 462125 213273
rect 475278 213404 475422 213408
rect 475278 213268 475282 213404
rect 475282 213268 475418 213404
rect 475418 213268 475422 213404
rect 475278 213264 475422 213268
rect 487626 213378 487770 213382
rect 487626 213242 487630 213378
rect 487630 213242 487766 213378
rect 487766 213242 487770 213378
rect 487626 213238 487770 213242
rect 534929 213154 535313 213538
rect 569529 213155 569913 213539
rect 86957 212762 87101 212766
rect 86957 212626 86961 212762
rect 86961 212626 87097 212762
rect 87097 212626 87101 212762
rect 86957 212622 87101 212626
rect 89719 212731 89863 212735
rect 89719 212595 89723 212731
rect 89723 212595 89859 212731
rect 89859 212595 89863 212731
rect 89719 212591 89863 212595
rect 99302 212711 99446 212715
rect 99302 212575 99306 212711
rect 99306 212575 99442 212711
rect 99442 212575 99446 212711
rect 99302 212571 99446 212575
rect 102075 212736 102219 212740
rect 102075 212600 102079 212736
rect 102079 212600 102215 212736
rect 102215 212600 102219 212736
rect 102075 212596 102219 212600
rect 112262 212746 112406 212750
rect 112262 212610 112266 212746
rect 112266 212610 112402 212746
rect 112402 212610 112406 212746
rect 112262 212606 112406 212610
rect 115029 212771 115173 212775
rect 115029 212635 115033 212771
rect 115033 212635 115169 212771
rect 115169 212635 115173 212771
rect 115029 212631 115173 212635
rect 124601 212736 124745 212740
rect 124601 212600 124605 212736
rect 124605 212600 124741 212736
rect 124741 212600 124745 212736
rect 124601 212596 124745 212600
rect 127374 212727 127518 212731
rect 127374 212591 127378 212727
rect 127378 212591 127514 212727
rect 127514 212591 127518 212727
rect 127374 212587 127518 212591
rect 137917 212723 138061 212727
rect 137917 212587 137921 212723
rect 137921 212587 138057 212723
rect 138057 212587 138061 212723
rect 137917 212583 138061 212587
rect 140679 212743 140823 212747
rect 140679 212607 140683 212743
rect 140683 212607 140819 212743
rect 140819 212607 140823 212743
rect 140679 212603 140823 212607
rect 150259 212684 150403 212688
rect 150259 212548 150263 212684
rect 150263 212548 150399 212684
rect 150399 212548 150403 212684
rect 150259 212544 150403 212548
rect 153017 212700 153161 212704
rect 153017 212564 153021 212700
rect 153021 212564 153157 212700
rect 153157 212564 153161 212700
rect 153017 212560 153161 212564
rect 163559 212701 163703 212705
rect 163559 212565 163563 212701
rect 163563 212565 163699 212701
rect 163699 212565 163703 212701
rect 163559 212561 163703 212565
rect 166330 212689 166474 212693
rect 166330 212553 166334 212689
rect 166334 212553 166470 212689
rect 166470 212553 166474 212689
rect 166330 212549 166474 212553
rect 175909 212708 176053 212712
rect 175909 212572 175913 212708
rect 175913 212572 176049 212708
rect 176049 212572 176053 212708
rect 175909 212568 176053 212572
rect 178670 212689 178814 212693
rect 178670 212553 178674 212689
rect 178674 212553 178810 212689
rect 178810 212553 178814 212689
rect 178670 212549 178814 212553
rect 189213 212715 189357 212719
rect 189213 212579 189217 212715
rect 189217 212579 189353 212715
rect 189353 212579 189357 212715
rect 189213 212575 189357 212579
rect 191980 212715 192124 212719
rect 191980 212579 191984 212715
rect 191984 212579 192120 212715
rect 192120 212579 192124 212715
rect 191980 212575 192124 212579
rect 201554 212725 201698 212729
rect 201554 212589 201558 212725
rect 201558 212589 201694 212725
rect 201694 212589 201698 212725
rect 201554 212585 201698 212589
rect 204320 212703 204464 212707
rect 204320 212567 204324 212703
rect 204324 212567 204460 212703
rect 204460 212567 204464 212703
rect 204320 212563 204464 212567
rect 214862 212745 215006 212749
rect 214862 212609 214866 212745
rect 214866 212609 215002 212745
rect 215002 212609 215006 212745
rect 214862 212605 215006 212609
rect 217626 212741 217770 212745
rect 217626 212605 217630 212741
rect 217630 212605 217766 212741
rect 217766 212605 217770 212741
rect 217626 212601 217770 212605
rect 227213 212734 227357 212738
rect 227213 212598 227217 212734
rect 227217 212598 227353 212734
rect 227353 212598 227357 212734
rect 227213 212594 227357 212598
rect 229972 212712 230116 212716
rect 229972 212576 229976 212712
rect 229976 212576 230112 212712
rect 230112 212576 230116 212712
rect 229972 212572 230116 212576
rect 240514 212733 240658 212737
rect 240514 212597 240518 212733
rect 240518 212597 240654 212733
rect 240654 212597 240658 212733
rect 240514 212593 240658 212597
rect 243275 212742 243419 212746
rect 243275 212606 243279 212742
rect 243279 212606 243415 212742
rect 243415 212606 243419 212742
rect 243275 212602 243419 212606
rect 252860 212723 253004 212727
rect 252860 212587 252864 212723
rect 252864 212587 253000 212723
rect 253000 212587 253004 212723
rect 252860 212583 253004 212587
rect 255620 212723 255764 212727
rect 255620 212587 255624 212723
rect 255624 212587 255760 212723
rect 255760 212587 255764 212723
rect 255620 212583 255764 212587
rect 266161 212639 266305 212643
rect 266161 212503 266165 212639
rect 266165 212503 266301 212639
rect 266301 212503 266305 212639
rect 266161 212499 266305 212503
rect 268928 212673 269072 212677
rect 268928 212537 268932 212673
rect 268932 212537 269068 212673
rect 269068 212537 269072 212673
rect 268928 212533 269072 212537
rect 278505 212704 278649 212708
rect 278505 212568 278509 212704
rect 278509 212568 278645 212704
rect 278645 212568 278649 212704
rect 278505 212564 278649 212568
rect 281273 212714 281417 212718
rect 281273 212578 281277 212714
rect 281277 212578 281413 212714
rect 281413 212578 281417 212714
rect 281273 212574 281417 212578
rect 291813 212648 291957 212652
rect 291813 212512 291817 212648
rect 291817 212512 291953 212648
rect 291953 212512 291957 212648
rect 291813 212508 291957 212512
rect 294576 212669 294720 212673
rect 294576 212533 294580 212669
rect 294580 212533 294716 212669
rect 294716 212533 294720 212669
rect 294576 212529 294720 212533
rect 304165 212689 304309 212693
rect 304165 212553 304169 212689
rect 304169 212553 304305 212689
rect 304305 212553 304309 212689
rect 304165 212549 304309 212553
rect 306929 212684 307073 212688
rect 306929 212548 306933 212684
rect 306933 212548 307069 212684
rect 307069 212548 307073 212684
rect 306929 212544 307073 212548
rect 317468 212704 317612 212708
rect 317468 212568 317472 212704
rect 317472 212568 317608 212704
rect 317608 212568 317612 212704
rect 317468 212564 317612 212568
rect 320226 212704 320370 212708
rect 320226 212568 320230 212704
rect 320230 212568 320366 212704
rect 320366 212568 320370 212704
rect 320226 212564 320370 212568
rect 329809 212731 329953 212735
rect 329809 212595 329813 212731
rect 329813 212595 329949 212731
rect 329949 212595 329953 212731
rect 329809 212591 329953 212595
rect 332572 212766 332716 212770
rect 332572 212630 332576 212766
rect 332576 212630 332712 212766
rect 332712 212630 332716 212766
rect 332572 212626 332716 212630
rect 343115 212702 343259 212706
rect 343115 212566 343119 212702
rect 343119 212566 343255 212702
rect 343255 212566 343259 212702
rect 343115 212562 343259 212566
rect 345877 212707 346021 212711
rect 345877 212571 345881 212707
rect 345881 212571 346017 212707
rect 346017 212571 346021 212707
rect 345877 212567 346021 212571
rect 355456 212698 355600 212702
rect 355456 212562 355460 212698
rect 355460 212562 355596 212698
rect 355596 212562 355600 212698
rect 355456 212558 355600 212562
rect 358222 212717 358366 212721
rect 358222 212581 358226 212717
rect 358226 212581 358362 212717
rect 358362 212581 358366 212717
rect 358222 212577 358366 212581
rect 368765 212684 368909 212688
rect 368765 212548 368769 212684
rect 368769 212548 368905 212684
rect 368905 212548 368909 212684
rect 368765 212544 368909 212548
rect 371527 212708 371671 212712
rect 371527 212572 371531 212708
rect 371531 212572 371667 212708
rect 371667 212572 371671 212708
rect 371527 212568 371671 212572
rect 381109 212731 381253 212735
rect 381109 212595 381113 212731
rect 381113 212595 381249 212731
rect 381249 212595 381253 212731
rect 381109 212591 381253 212595
rect 383874 212750 384018 212754
rect 383874 212614 383878 212750
rect 383878 212614 384014 212750
rect 384014 212614 384018 212750
rect 383874 212610 384018 212614
rect 394416 212695 394560 212699
rect 394416 212559 394420 212695
rect 394420 212559 394556 212695
rect 394556 212559 394560 212695
rect 394416 212555 394560 212559
rect 397177 212745 397321 212749
rect 397177 212609 397181 212745
rect 397181 212609 397317 212745
rect 397317 212609 397321 212745
rect 397177 212605 397321 212609
rect 406755 212711 406899 212715
rect 406755 212575 406759 212711
rect 406759 212575 406895 212711
rect 406895 212575 406899 212711
rect 406755 212571 406899 212575
rect 409524 212731 409668 212735
rect 409524 212595 409528 212731
rect 409528 212595 409664 212731
rect 409664 212595 409668 212731
rect 409524 212591 409668 212595
rect 420065 212736 420209 212740
rect 420065 212600 420069 212736
rect 420069 212600 420205 212736
rect 420205 212600 420209 212736
rect 420065 212596 420209 212600
rect 422828 212754 422972 212758
rect 422828 212618 422832 212754
rect 422832 212618 422968 212754
rect 422968 212618 422972 212754
rect 422828 212614 422972 212618
rect 432414 212751 432558 212755
rect 432414 212615 432418 212751
rect 432418 212615 432554 212751
rect 432554 212615 432558 212751
rect 432414 212611 432558 212615
rect 435173 212723 435317 212727
rect 435173 212587 435177 212723
rect 435177 212587 435313 212723
rect 435313 212587 435317 212723
rect 435173 212583 435317 212587
rect 445709 212668 445853 212672
rect 445709 212532 445713 212668
rect 445713 212532 445849 212668
rect 445849 212532 445853 212668
rect 445709 212528 445853 212532
rect 448477 212722 448621 212726
rect 448477 212586 448481 212722
rect 448481 212586 448617 212722
rect 448617 212586 448621 212722
rect 448477 212582 448621 212586
rect 458059 212683 458203 212687
rect 458059 212547 458063 212683
rect 458063 212547 458199 212683
rect 458199 212547 458203 212683
rect 458059 212543 458203 212547
rect 460821 212715 460965 212719
rect 460821 212579 460825 212715
rect 460825 212579 460961 212715
rect 460961 212579 460965 212715
rect 460821 212575 460965 212579
rect 471356 212637 471500 212641
rect 471356 212501 471360 212637
rect 471360 212501 471496 212637
rect 471496 212501 471500 212637
rect 471356 212497 471500 212501
rect 474128 212691 474272 212695
rect 474128 212555 474132 212691
rect 474132 212555 474268 212691
rect 474268 212555 474272 212691
rect 474128 212551 474272 212555
rect 483712 212649 483856 212653
rect 483712 212513 483716 212649
rect 483716 212513 483852 212649
rect 483852 212513 483856 212649
rect 483712 212509 483856 212513
rect 486475 212719 486619 212723
rect 486475 212583 486479 212719
rect 486479 212583 486615 212719
rect 486615 212583 486619 212719
rect 486475 212579 486619 212583
rect 570135 144511 570519 144895
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 522682 688496 523482 688504
rect 512517 688454 513317 688462
rect 172220 688024 172620 688032
rect 95437 687801 95837 687809
rect 95437 687417 95445 687801
rect 95829 687417 95837 687801
rect 172220 687640 172228 688024
rect 172612 687640 172620 688024
rect 454201 687699 454601 687707
rect 172220 687632 172620 687640
rect 223339 687659 223739 687667
rect 95437 687409 95837 687417
rect 120762 687615 121162 687623
rect 120762 687231 120770 687615
rect 121154 687231 121162 687615
rect 216358 687584 216758 687592
rect 120762 687223 121162 687231
rect 146419 687493 146819 687501
rect 146419 687109 146427 687493
rect 146811 687109 146819 687493
rect 216358 687200 216366 687584
rect 216750 687200 216758 687584
rect 223339 687275 223347 687659
rect 223731 687275 223739 687659
rect 412441 687640 412841 687648
rect 300303 687614 300703 687622
rect 274678 687578 275078 687586
rect 223339 687267 223739 687275
rect 249009 687562 249409 687570
rect 216358 687192 216758 687200
rect 249009 687178 249017 687562
rect 249401 687178 249409 687562
rect 274678 687194 274686 687578
rect 275070 687194 275078 687578
rect 300303 687230 300311 687614
rect 300695 687230 300703 687614
rect 300303 687222 300703 687230
rect 325939 687579 326339 687587
rect 274678 687186 275078 687194
rect 325939 687195 325947 687579
rect 326331 687195 326339 687579
rect 325939 687187 326339 687195
rect 351604 687561 352004 687569
rect 249009 687170 249409 687178
rect 351604 687177 351612 687561
rect 351996 687177 352004 687561
rect 351604 687169 352004 687177
rect 377265 687523 377665 687531
rect 377265 687139 377273 687523
rect 377657 687139 377665 687523
rect 412441 687256 412449 687640
rect 412833 687256 412841 687640
rect 412441 687248 412841 687256
rect 428567 687630 428967 687638
rect 428567 687246 428575 687630
rect 428959 687246 428967 687630
rect 454201 687315 454209 687699
rect 454593 687315 454601 687699
rect 454201 687307 454601 687315
rect 479850 687705 480250 687713
rect 479850 687321 479858 687705
rect 480242 687321 480250 687705
rect 512517 687670 512525 688454
rect 513309 687670 513317 688454
rect 522682 687712 522690 688496
rect 523474 687712 523482 688496
rect 522682 687704 523482 687712
rect 512517 687662 513317 687670
rect 479850 687313 480250 687321
rect 428567 687238 428967 687246
rect 377265 687131 377665 687139
rect 146419 687101 146819 687109
rect 16246 678007 549815 680407
rect 10426 531016 10826 531024
rect 10426 530632 10434 531016
rect 10818 530632 10826 531016
rect 10426 530624 10826 530632
rect 9834 214911 10234 214919
rect 9834 214527 9842 214911
rect 10226 214527 10234 214911
rect 9834 214519 10234 214527
rect 16246 212880 18646 678007
rect 547415 621493 549815 678007
rect 560425 644576 566979 644980
rect 560425 639792 560582 644576
rect 566726 639792 566979 644576
rect 560425 634576 566979 639792
rect 560425 629792 560582 634576
rect 566726 629792 566979 634576
rect 560425 621493 566979 629792
rect 547415 619093 566979 621493
rect 37851 542711 38251 542719
rect 37851 542327 37859 542711
rect 38243 542327 38251 542711
rect 37851 542319 38251 542327
rect 75600 438027 76400 438200
rect 75600 437883 76152 438027
rect 76296 437883 76400 438027
rect 75600 435271 76400 437883
rect 75600 435127 76169 435271
rect 76313 435127 76400 435271
rect 75600 424687 76400 435127
rect 76998 434169 77398 434251
rect 76998 433933 77080 434169
rect 77316 433933 77398 434169
rect 76998 433851 77398 433933
rect 78895 433228 79295 433310
rect 78895 432992 78977 433228
rect 79213 432992 79295 433228
rect 78895 432910 79295 432992
rect 75600 424543 76179 424687
rect 76323 424543 76400 424687
rect 75600 421921 76400 424543
rect 75600 421777 76194 421921
rect 76338 421777 76400 421921
rect 75600 411343 76400 421777
rect 76998 420824 77398 420906
rect 76998 420588 77080 420824
rect 77316 420588 77398 420824
rect 76998 420506 77398 420588
rect 78896 419869 79296 419951
rect 78896 419633 78978 419869
rect 79214 419633 79296 419869
rect 78896 419551 79296 419633
rect 75600 411199 76163 411343
rect 76307 411199 76400 411343
rect 75600 408576 76400 411199
rect 75600 408432 76194 408576
rect 76338 408432 76400 408576
rect 75600 397988 76400 408432
rect 76998 407470 77398 407552
rect 76998 407234 77080 407470
rect 77316 407234 77398 407470
rect 76998 407152 77398 407234
rect 78897 406530 79297 406612
rect 78897 406294 78979 406530
rect 79215 406294 79297 406530
rect 78897 406212 79297 406294
rect 75600 397844 76176 397988
rect 76320 397844 76400 397988
rect 75600 395234 76400 397844
rect 75600 395090 76181 395234
rect 76325 395090 76400 395234
rect 75600 384648 76400 395090
rect 76998 394147 77398 394229
rect 76998 393911 77080 394147
rect 77316 393911 77398 394147
rect 76998 393829 77398 393911
rect 78896 393195 79296 393277
rect 78896 392959 78978 393195
rect 79214 392959 79296 393195
rect 78896 392877 79296 392959
rect 75600 384504 76151 384648
rect 76295 384504 76400 384648
rect 75600 381886 76400 384504
rect 75600 381742 76156 381886
rect 76300 381742 76400 381886
rect 75600 371306 76400 381742
rect 76998 380781 77398 380863
rect 76998 380545 77080 380781
rect 77316 380545 77398 380781
rect 76998 380463 77398 380545
rect 78896 379842 79296 379924
rect 78896 379606 78978 379842
rect 79214 379606 79296 379842
rect 78896 379524 79296 379606
rect 75600 371162 76171 371306
rect 76315 371162 76400 371306
rect 75600 368545 76400 371162
rect 75600 368401 76174 368545
rect 76318 368401 76400 368545
rect 75600 357957 76400 368401
rect 76998 367427 77398 367509
rect 76998 367191 77080 367427
rect 77316 367191 77398 367427
rect 76998 367109 77398 367191
rect 78898 366486 79298 366568
rect 78898 366250 78980 366486
rect 79216 366250 79298 366486
rect 78898 366168 79298 366250
rect 75600 357813 76161 357957
rect 76305 357813 76400 357957
rect 75600 355200 76400 357813
rect 75600 355056 76181 355200
rect 76325 355056 76400 355200
rect 75600 344612 76400 355056
rect 76998 354090 77398 354172
rect 76998 353854 77080 354090
rect 77316 354041 77398 354090
rect 77317 353897 77398 354041
rect 77316 353854 77398 353897
rect 76998 353772 77398 353854
rect 78896 353158 79296 353240
rect 78896 352922 78978 353158
rect 79214 352922 79296 353158
rect 78896 352840 79296 352922
rect 75600 344468 76128 344612
rect 76272 344468 76400 344612
rect 75600 341850 76400 344468
rect 75600 341706 76151 341850
rect 76295 341706 76400 341850
rect 75600 331268 76400 341706
rect 77000 340741 77400 340823
rect 77000 340505 77082 340741
rect 77318 340505 77400 340741
rect 77000 340423 77400 340505
rect 78898 339813 79298 339895
rect 78898 339577 78980 339813
rect 79216 339577 79298 339813
rect 78898 339495 79298 339577
rect 75600 331124 76171 331268
rect 76315 331124 76400 331268
rect 75600 328510 76400 331124
rect 75600 328366 76175 328510
rect 76319 328366 76400 328510
rect 75600 317916 76400 328366
rect 76999 327376 77399 327458
rect 76999 327140 77081 327376
rect 77317 327140 77399 327376
rect 76999 327058 77399 327140
rect 78894 326461 79294 326543
rect 78894 326225 78976 326461
rect 79212 326225 79294 326461
rect 78894 326143 79294 326225
rect 75600 317772 76183 317916
rect 76327 317772 76400 317916
rect 75600 315165 76400 317772
rect 75600 315021 76171 315165
rect 76315 315021 76400 315165
rect 75600 304575 76400 315021
rect 76998 314049 77398 314131
rect 76998 313813 77080 314049
rect 77316 313813 77398 314049
rect 76998 313731 77398 313813
rect 78897 313094 79297 313176
rect 78897 312858 78979 313094
rect 79215 312858 79297 313094
rect 78897 312776 79297 312858
rect 75600 304431 76166 304575
rect 76310 304431 76400 304575
rect 75600 301818 76400 304431
rect 75600 301674 76181 301818
rect 76325 301674 76400 301818
rect 75600 291235 76400 301674
rect 76998 300693 77398 300775
rect 76998 300457 77080 300693
rect 77316 300457 77398 300693
rect 76998 300375 77398 300457
rect 78895 299773 79295 299855
rect 78895 299537 78977 299773
rect 79213 299537 79295 299773
rect 78895 299455 79295 299537
rect 75600 291091 76166 291235
rect 76310 291091 76400 291235
rect 75600 288482 76400 291091
rect 75600 288338 76156 288482
rect 76300 288338 76400 288482
rect 75600 277901 76400 288338
rect 76998 287354 77398 287436
rect 76998 287118 77080 287354
rect 77316 287118 77398 287354
rect 76998 287036 77398 287118
rect 78894 286412 79294 286494
rect 78894 286176 78976 286412
rect 79212 286176 79294 286412
rect 78894 286094 79294 286176
rect 75600 277757 76174 277901
rect 76318 277757 76400 277901
rect 75600 275123 76400 277757
rect 75600 274979 76174 275123
rect 76318 274979 76400 275123
rect 75600 264544 76400 274979
rect 76999 274020 77399 274102
rect 76999 273784 77081 274020
rect 77317 273784 77399 274020
rect 76999 273702 77399 273784
rect 78897 273072 79297 273154
rect 78897 272836 78979 273072
rect 79215 272836 79297 273072
rect 78897 272754 79297 272836
rect 75600 264400 76185 264544
rect 76329 264400 76400 264544
rect 75600 261785 76400 264400
rect 75600 261641 76197 261785
rect 76341 261641 76400 261785
rect 75600 251195 76400 261641
rect 76999 260672 77399 260754
rect 76999 260436 77081 260672
rect 77317 260436 77399 260672
rect 76999 260354 77399 260436
rect 78896 259728 79296 259810
rect 78896 259492 78978 259728
rect 79214 259492 79296 259728
rect 78896 259410 79296 259492
rect 75600 251051 76182 251195
rect 76326 251051 76400 251195
rect 75600 248436 76400 251051
rect 75600 248292 76180 248436
rect 76324 248292 76400 248436
rect 75600 237850 76400 248292
rect 76998 247322 77398 247404
rect 76998 247086 77080 247322
rect 77316 247086 77398 247322
rect 76998 247004 77398 247086
rect 78896 246374 79296 246456
rect 78896 246138 78978 246374
rect 79214 246138 79296 246374
rect 78896 246056 79296 246138
rect 75600 237822 76401 237850
rect 75600 237678 76229 237822
rect 76373 237678 76401 237822
rect 75600 237650 76401 237678
rect 75600 235054 76400 237650
rect 75600 234910 76227 235054
rect 76371 234910 76400 235054
rect 75600 212880 76400 234910
rect 76997 233955 77397 234037
rect 76997 233719 77079 233955
rect 77315 233719 77397 233955
rect 76997 233637 77397 233719
rect 539186 233284 540786 233292
rect 78881 232990 79281 233072
rect 78881 232754 78963 232990
rect 79199 232754 79281 232990
rect 78881 232672 79281 232754
rect 539186 231700 539194 233284
rect 540778 231700 540786 233284
rect 539186 231692 540786 231700
rect 91696 215254 92096 215336
rect 91696 215018 91778 215254
rect 92014 215018 92096 215254
rect 91696 214936 92096 215018
rect 104041 215259 104441 215341
rect 104041 215023 104123 215259
rect 104359 215023 104441 215259
rect 104041 214941 104441 215023
rect 117001 215245 117401 215327
rect 117001 215009 117083 215245
rect 117319 215009 117401 215245
rect 117001 214927 117401 215009
rect 129354 215255 129754 215337
rect 129354 215019 129436 215255
rect 129672 215019 129754 215255
rect 129354 214937 129754 215019
rect 142659 215254 143059 215336
rect 142659 215018 142741 215254
rect 142977 215018 143059 215254
rect 142659 214936 143059 215018
rect 155003 215256 155403 215338
rect 155003 215020 155085 215256
rect 155321 215020 155403 215256
rect 155003 214938 155403 215020
rect 168306 215258 168706 215340
rect 168306 215022 168388 215258
rect 168624 215022 168706 215258
rect 168306 214940 168706 215022
rect 180652 215259 181052 215341
rect 180652 215023 180734 215259
rect 180970 215023 181052 215259
rect 180652 214941 181052 215023
rect 193943 215265 194343 215347
rect 193943 215029 194025 215265
rect 194261 215029 194343 215265
rect 193943 214947 194343 215029
rect 206288 215258 206688 215340
rect 206288 215022 206370 215258
rect 206606 215022 206688 215258
rect 206288 214940 206688 215022
rect 219598 215256 219998 215338
rect 219598 215020 219680 215256
rect 219916 215020 219998 215256
rect 219598 214938 219998 215020
rect 231942 215257 232342 215331
rect 231942 215249 232074 215257
rect 232218 215249 232342 215257
rect 231942 215013 232024 215249
rect 232260 215013 232342 215249
rect 231942 214931 232342 215013
rect 245244 215264 245644 215346
rect 245244 215028 245326 215264
rect 245562 215028 245644 215264
rect 245244 214946 245644 215028
rect 257586 215272 257986 215340
rect 257586 215258 257723 215272
rect 257867 215258 257986 215272
rect 257586 215022 257668 215258
rect 257904 215022 257986 215258
rect 257586 214940 257986 215022
rect 270905 215258 271305 215340
rect 270905 215022 270987 215258
rect 271223 215022 271305 215258
rect 270905 214940 271305 215022
rect 283237 215261 283637 215343
rect 283237 215025 283319 215261
rect 283555 215025 283637 215261
rect 283237 214943 283637 215025
rect 296542 215254 296942 215336
rect 296542 215018 296624 215254
rect 296860 215018 296942 215254
rect 296542 214936 296942 215018
rect 308898 215258 309298 215340
rect 308898 215022 308980 215258
rect 309216 215022 309298 215258
rect 308898 214940 309298 215022
rect 322175 215245 322575 215327
rect 322175 215009 322257 215245
rect 322493 215009 322575 215245
rect 322175 214927 322575 215009
rect 334543 215256 334943 215338
rect 334543 215020 334625 215256
rect 334861 215020 334943 215256
rect 334543 214938 334943 215020
rect 347846 215263 348246 215345
rect 347846 215027 347928 215263
rect 348164 215027 348246 215263
rect 347846 214945 348246 215027
rect 360200 215256 360600 215338
rect 360200 215020 360282 215256
rect 360518 215020 360600 215256
rect 360200 214938 360600 215020
rect 373494 215249 373894 215331
rect 373494 215013 373576 215249
rect 373812 215013 373894 215249
rect 373494 214931 373894 215013
rect 385836 215259 386236 215341
rect 385836 215023 385918 215259
rect 386154 215023 386236 215259
rect 385836 214941 386236 215023
rect 399153 215256 399553 215338
rect 399153 215020 399235 215256
rect 399471 215020 399553 215256
rect 399153 214938 399553 215020
rect 411484 215259 411884 215341
rect 411484 215023 411566 215259
rect 411802 215023 411884 215259
rect 411484 214941 411884 215023
rect 424803 215258 425203 215340
rect 424803 215022 424885 215258
rect 425121 215022 425203 215258
rect 424803 214940 425203 215022
rect 437143 215258 437543 215340
rect 437143 215022 437225 215258
rect 437461 215022 437543 215258
rect 437143 214940 437543 215022
rect 450439 215258 450839 215340
rect 450439 215022 450521 215258
rect 450757 215022 450839 215258
rect 450439 214940 450839 215022
rect 462803 215261 463203 215343
rect 462803 215025 462885 215261
rect 463121 215025 463203 215261
rect 462803 214943 463203 215025
rect 476105 215259 476505 215341
rect 476105 215023 476187 215259
rect 476423 215023 476505 215259
rect 476105 214941 476505 215023
rect 488456 215259 488856 215341
rect 488456 215023 488538 215259
rect 488774 215023 488856 215259
rect 488456 214941 488856 215023
rect 90738 213466 91138 213548
rect 90738 213230 90820 213466
rect 91056 213230 91138 213466
rect 90738 213148 91138 213230
rect 103099 213461 103499 213543
rect 103099 213225 103181 213461
rect 103417 213225 103499 213461
rect 103099 213143 103499 213225
rect 116063 213470 116463 213552
rect 116063 213234 116145 213470
rect 116381 213234 116463 213470
rect 116063 213152 116463 213234
rect 128396 213458 128796 213540
rect 128396 213222 128478 213458
rect 128714 213222 128796 213458
rect 128396 213140 128796 213222
rect 141701 213447 142101 213529
rect 141701 213211 141783 213447
rect 142019 213211 142101 213447
rect 141701 213201 141829 213211
rect 141973 213201 142101 213211
rect 141701 213129 142101 213201
rect 154044 213460 154444 213542
rect 154044 213224 154126 213460
rect 154362 213224 154444 213460
rect 154044 213142 154444 213224
rect 167350 213460 167750 213542
rect 167350 213224 167432 213460
rect 167668 213224 167750 213460
rect 167350 213142 167750 213224
rect 179709 213464 180109 213546
rect 179709 213228 179791 213464
rect 180027 213228 180109 213464
rect 179709 213146 180109 213228
rect 192987 213464 193387 213546
rect 192987 213228 193069 213464
rect 193305 213228 193387 213464
rect 192987 213146 193387 213228
rect 205346 213471 205746 213553
rect 205346 213235 205428 213471
rect 205664 213235 205746 213471
rect 205346 213153 205746 213235
rect 218648 213464 219048 213546
rect 218648 213228 218730 213464
rect 218966 213228 219048 213464
rect 218648 213146 219048 213228
rect 230992 213462 231392 213544
rect 230992 213226 231074 213462
rect 231310 213226 231392 213462
rect 230992 213144 231392 213226
rect 244286 213458 244686 213540
rect 244286 213222 244368 213458
rect 244604 213222 244686 213458
rect 244286 213140 244686 213222
rect 256653 213464 257053 213546
rect 256653 213228 256735 213464
rect 256971 213228 257053 213464
rect 256653 213146 257053 213228
rect 269959 213457 270359 213539
rect 269959 213221 270041 213457
rect 270277 213221 270359 213457
rect 269959 213139 270359 213221
rect 282285 213463 282685 213545
rect 282285 213227 282367 213463
rect 282603 213227 282685 213463
rect 282285 213223 282430 213227
rect 282574 213223 282685 213227
rect 282285 213145 282685 213223
rect 295596 213460 295996 213542
rect 295596 213224 295678 213460
rect 295914 213224 295996 213460
rect 295596 213142 295996 213224
rect 307944 213453 308344 213535
rect 307944 213217 308026 213453
rect 308262 213217 308344 213453
rect 307944 213196 308081 213217
rect 308225 213196 308344 213217
rect 307944 213135 308344 213196
rect 321251 213458 321651 213540
rect 321251 213222 321333 213458
rect 321569 213222 321651 213458
rect 321251 213140 321651 213222
rect 333606 213460 334006 213542
rect 333606 213224 333688 213460
rect 333924 213224 334006 213460
rect 333606 213212 333724 213224
rect 333868 213212 334006 213224
rect 333606 213142 334006 213212
rect 346888 213463 347288 213545
rect 346888 213227 346970 213463
rect 347206 213227 347288 213463
rect 346888 213145 347288 213227
rect 359228 213463 359628 213545
rect 359228 213227 359310 213463
rect 359546 213227 359628 213463
rect 359228 213145 359628 213227
rect 372557 213464 372957 213546
rect 372557 213228 372639 213464
rect 372875 213228 372957 213464
rect 372557 213146 372957 213228
rect 384900 213464 385300 213546
rect 384900 213228 384982 213464
rect 385218 213228 385300 213464
rect 384900 213146 385300 213228
rect 398190 213464 398590 213546
rect 398190 213228 398272 213464
rect 398508 213228 398590 213464
rect 398190 213146 398590 213228
rect 410539 213467 410939 213549
rect 410539 213231 410621 213467
rect 410857 213231 410939 213467
rect 410539 213149 410939 213231
rect 423859 213466 424259 213548
rect 423859 213230 423941 213466
rect 424177 213230 424259 213466
rect 423859 213148 424259 213230
rect 436200 213535 436600 213543
rect 436200 213151 436208 213535
rect 436592 213151 436600 213535
rect 436200 213143 436600 213151
rect 449509 213459 449909 213541
rect 449509 213223 449591 213459
rect 449827 213223 449909 213459
rect 449509 213141 449909 213223
rect 461861 213462 462261 213544
rect 461861 213226 461943 213462
rect 462179 213226 462261 213462
rect 461861 213144 462261 213226
rect 475141 213458 475541 213540
rect 475141 213222 475223 213458
rect 475459 213222 475541 213458
rect 475141 213140 475541 213222
rect 487497 213463 487897 213545
rect 487497 213227 487579 213463
rect 487815 213227 487897 213463
rect 487497 213145 487897 213227
rect 534921 213538 535321 213546
rect 534921 213154 534929 213538
rect 535313 213154 535321 213538
rect 534921 213146 535321 213154
rect 16246 212775 497417 212880
rect 16246 212766 115029 212775
rect 16246 212622 86957 212766
rect 87101 212750 115029 212766
rect 87101 212740 112262 212750
rect 87101 212735 102075 212740
rect 87101 212622 89719 212735
rect 16246 212591 89719 212622
rect 89863 212715 102075 212735
rect 89863 212591 99302 212715
rect 16246 212571 99302 212591
rect 99446 212596 102075 212715
rect 102219 212606 112262 212740
rect 112406 212631 115029 212750
rect 115173 212770 497417 212775
rect 115173 212749 332572 212770
rect 115173 212747 214862 212749
rect 115173 212740 140679 212747
rect 115173 212631 124601 212740
rect 112406 212606 124601 212631
rect 102219 212596 124601 212606
rect 124745 212731 140679 212740
rect 124745 212596 127374 212731
rect 99446 212587 127374 212596
rect 127518 212727 140679 212731
rect 127518 212587 137917 212727
rect 99446 212583 137917 212587
rect 138061 212603 140679 212727
rect 140823 212729 214862 212747
rect 140823 212719 201554 212729
rect 140823 212712 189213 212719
rect 140823 212705 175909 212712
rect 140823 212704 163559 212705
rect 140823 212688 153017 212704
rect 140823 212603 150259 212688
rect 138061 212583 150259 212603
rect 99446 212571 150259 212583
rect 16246 212544 150259 212571
rect 150403 212560 153017 212688
rect 153161 212561 163559 212704
rect 163703 212693 175909 212705
rect 163703 212561 166330 212693
rect 153161 212560 166330 212561
rect 150403 212549 166330 212560
rect 166474 212568 175909 212693
rect 176053 212693 189213 212712
rect 176053 212568 178670 212693
rect 166474 212549 178670 212568
rect 178814 212575 189213 212693
rect 189357 212575 191980 212719
rect 192124 212585 201554 212719
rect 201698 212707 214862 212729
rect 201698 212585 204320 212707
rect 192124 212575 204320 212585
rect 178814 212563 204320 212575
rect 204464 212605 214862 212707
rect 215006 212746 332572 212749
rect 215006 212745 243275 212746
rect 215006 212605 217626 212745
rect 204464 212601 217626 212605
rect 217770 212738 243275 212745
rect 217770 212601 227213 212738
rect 204464 212594 227213 212601
rect 227357 212737 243275 212738
rect 227357 212716 240514 212737
rect 227357 212594 229972 212716
rect 204464 212572 229972 212594
rect 230116 212593 240514 212716
rect 240658 212602 243275 212737
rect 243419 212735 332572 212746
rect 243419 212727 329809 212735
rect 243419 212602 252860 212727
rect 240658 212593 252860 212602
rect 230116 212583 252860 212593
rect 253004 212583 255620 212727
rect 255764 212718 329809 212727
rect 255764 212708 281273 212718
rect 255764 212677 278505 212708
rect 255764 212643 268928 212677
rect 255764 212583 266161 212643
rect 230116 212572 266161 212583
rect 204464 212563 266161 212572
rect 178814 212549 266161 212563
rect 150403 212544 266161 212549
rect 16246 212499 266161 212544
rect 266305 212533 268928 212643
rect 269072 212564 278505 212677
rect 278649 212574 281273 212708
rect 281417 212708 329809 212718
rect 281417 212693 317468 212708
rect 281417 212673 304165 212693
rect 281417 212652 294576 212673
rect 281417 212574 291813 212652
rect 278649 212564 291813 212574
rect 269072 212533 291813 212564
rect 266305 212508 291813 212533
rect 291957 212529 294576 212652
rect 294720 212549 304165 212673
rect 304309 212688 317468 212693
rect 304309 212549 306929 212688
rect 294720 212544 306929 212549
rect 307073 212564 317468 212688
rect 317612 212564 320226 212708
rect 320370 212591 329809 212708
rect 329953 212626 332572 212735
rect 332716 212758 497417 212770
rect 332716 212754 422828 212758
rect 332716 212735 383874 212754
rect 332716 212721 381109 212735
rect 332716 212711 358222 212721
rect 332716 212706 345877 212711
rect 332716 212626 343115 212706
rect 329953 212591 343115 212626
rect 320370 212564 343115 212591
rect 307073 212562 343115 212564
rect 343259 212567 345877 212706
rect 346021 212702 358222 212711
rect 346021 212567 355456 212702
rect 343259 212562 355456 212567
rect 307073 212558 355456 212562
rect 355600 212577 358222 212702
rect 358366 212712 381109 212721
rect 358366 212688 371527 212712
rect 358366 212577 368765 212688
rect 355600 212558 368765 212577
rect 307073 212544 368765 212558
rect 368909 212568 371527 212688
rect 371671 212591 381109 212712
rect 381253 212610 383874 212735
rect 384018 212749 422828 212754
rect 384018 212699 397177 212749
rect 384018 212610 394416 212699
rect 381253 212591 394416 212610
rect 371671 212568 394416 212591
rect 368909 212555 394416 212568
rect 394560 212605 397177 212699
rect 397321 212740 422828 212749
rect 397321 212735 420065 212740
rect 397321 212715 409524 212735
rect 397321 212605 406755 212715
rect 394560 212571 406755 212605
rect 406899 212591 409524 212715
rect 409668 212596 420065 212735
rect 420209 212614 422828 212740
rect 422972 212755 497417 212758
rect 422972 212614 432414 212755
rect 420209 212611 432414 212614
rect 432558 212727 497417 212755
rect 432558 212611 435173 212727
rect 420209 212596 435173 212611
rect 409668 212591 435173 212596
rect 406899 212583 435173 212591
rect 435317 212726 497417 212727
rect 435317 212672 448477 212726
rect 435317 212583 445709 212672
rect 406899 212571 445709 212583
rect 394560 212555 445709 212571
rect 368909 212544 445709 212555
rect 294720 212529 445709 212544
rect 291957 212528 445709 212529
rect 445853 212582 448477 212672
rect 448621 212723 497417 212726
rect 448621 212719 486475 212723
rect 448621 212687 460821 212719
rect 448621 212582 458059 212687
rect 445853 212543 458059 212582
rect 458203 212575 460821 212687
rect 460965 212695 486475 212719
rect 460965 212641 474128 212695
rect 460965 212575 471356 212641
rect 458203 212543 471356 212575
rect 445853 212528 471356 212543
rect 291957 212508 471356 212528
rect 266305 212499 471356 212508
rect 16246 212497 471356 212499
rect 471500 212551 474128 212641
rect 474272 212653 486475 212695
rect 474272 212551 483712 212653
rect 471500 212509 483712 212551
rect 483856 212579 486475 212653
rect 486619 212579 497417 212723
rect 483856 212509 497417 212579
rect 471500 212497 497417 212509
rect 16246 212080 497417 212497
rect 16246 29052 18646 212080
rect 547415 29052 549815 619093
rect 560425 613756 566979 619093
rect 556059 555354 562613 595202
rect 556059 550570 556255 555354
rect 562319 550570 562613 555354
rect 556059 545354 562613 550570
rect 556059 540570 556255 545354
rect 562319 540570 562613 545354
rect 556059 540155 562613 540570
rect 569780 531017 570180 531025
rect 569780 530633 569788 531017
rect 570172 530633 570180 531017
rect 569780 530625 570180 530633
rect 569521 213539 569921 213547
rect 569521 213155 569529 213539
rect 569913 213155 569921 213539
rect 569521 213147 569921 213155
rect 570127 144895 570527 144903
rect 570127 144511 570135 144895
rect 570519 144511 570527 144895
rect 570127 144503 570527 144511
rect 16246 26652 549815 29052
<< via4 >>
rect 95519 687491 95755 687727
rect 172302 687714 172538 687950
rect 120844 687305 121080 687541
rect 146501 687183 146737 687419
rect 216440 687274 216676 687510
rect 223421 687349 223657 687585
rect 249091 687252 249327 687488
rect 274760 687268 274996 687504
rect 300385 687304 300621 687540
rect 326021 687269 326257 687505
rect 351686 687251 351922 687487
rect 377347 687213 377583 687449
rect 412523 687330 412759 687566
rect 428649 687320 428885 687556
rect 454283 687389 454519 687625
rect 479932 687395 480168 687631
rect 512639 687784 513195 688340
rect 522804 687826 523360 688382
rect 10508 530706 10744 530942
rect 9916 214601 10152 214837
rect 37933 542401 38169 542637
rect 77080 434115 77316 434169
rect 77080 433971 77100 434115
rect 77100 433971 77244 434115
rect 77244 433971 77316 434115
rect 77080 433933 77316 433971
rect 78977 433167 79213 433228
rect 78977 433023 79031 433167
rect 79031 433023 79175 433167
rect 79175 433023 79213 433167
rect 78977 432992 79213 433023
rect 77080 420763 77316 420824
rect 77080 420619 77133 420763
rect 77133 420619 77277 420763
rect 77277 420619 77316 420763
rect 77080 420588 77316 420619
rect 78978 419820 79214 419869
rect 78978 419676 79022 419820
rect 79022 419676 79166 419820
rect 79166 419676 79214 419820
rect 78978 419633 79214 419676
rect 77080 407423 77316 407470
rect 77080 407279 77121 407423
rect 77121 407279 77265 407423
rect 77265 407279 77316 407423
rect 77080 407234 77316 407279
rect 78979 406475 79215 406530
rect 78979 406331 79006 406475
rect 79006 406331 79150 406475
rect 79150 406331 79215 406475
rect 78979 406294 79215 406331
rect 77080 394074 77316 394147
rect 77080 393930 77133 394074
rect 77133 393930 77277 394074
rect 77277 393930 77316 394074
rect 77080 393911 77316 393930
rect 78978 393135 79214 393195
rect 78978 392991 79031 393135
rect 79031 392991 79175 393135
rect 79175 392991 79214 393135
rect 78978 392959 79214 392991
rect 77080 380730 77316 380781
rect 77080 380586 77121 380730
rect 77121 380586 77265 380730
rect 77265 380586 77316 380730
rect 77080 380545 77316 380586
rect 78978 379788 79214 379842
rect 78978 379644 78997 379788
rect 78997 379644 79141 379788
rect 79141 379644 79214 379788
rect 78978 379606 79214 379644
rect 77080 367385 77316 367427
rect 77080 367241 77083 367385
rect 77083 367241 77227 367385
rect 77227 367241 77316 367385
rect 77080 367191 77316 367241
rect 78980 366439 79216 366486
rect 78980 366295 79016 366439
rect 79016 366295 79160 366439
rect 79160 366295 79216 366439
rect 78980 366250 79216 366295
rect 77080 354041 77316 354090
rect 77080 353897 77173 354041
rect 77173 353897 77316 354041
rect 77080 353854 77316 353897
rect 78978 353099 79214 353158
rect 78978 352955 79020 353099
rect 79020 352955 79164 353099
rect 79164 352955 79214 353099
rect 78978 352922 79214 352955
rect 77082 340699 77318 340741
rect 77082 340555 77139 340699
rect 77139 340555 77283 340699
rect 77283 340555 77318 340699
rect 77082 340505 77318 340555
rect 78980 339750 79216 339813
rect 78980 339606 79027 339750
rect 79027 339606 79171 339750
rect 79171 339606 79216 339750
rect 78980 339577 79216 339606
rect 77081 327356 77317 327376
rect 77081 327212 77127 327356
rect 77127 327212 77271 327356
rect 77271 327212 77317 327356
rect 77081 327140 77317 327212
rect 78976 326402 79212 326461
rect 78976 326258 79039 326402
rect 79039 326258 79183 326402
rect 79183 326258 79212 326402
rect 78976 326225 79212 326258
rect 77080 314010 77316 314049
rect 77080 313866 77132 314010
rect 77132 313866 77276 314010
rect 77276 313866 77316 314010
rect 77080 313813 77316 313866
rect 78979 313064 79215 313094
rect 78979 312920 78998 313064
rect 78998 312920 79142 313064
rect 79142 312920 79215 313064
rect 78979 312858 79215 312920
rect 77080 300659 77316 300693
rect 77080 300515 77138 300659
rect 77138 300515 77282 300659
rect 77282 300515 77316 300659
rect 77080 300457 77316 300515
rect 78977 299713 79213 299773
rect 78977 299569 79011 299713
rect 79011 299569 79155 299713
rect 79155 299569 79213 299713
rect 78977 299537 79213 299569
rect 77080 287316 77316 287354
rect 77080 287172 77135 287316
rect 77135 287172 77279 287316
rect 77279 287172 77316 287316
rect 77080 287118 77316 287172
rect 78976 286370 79212 286412
rect 78976 286226 79009 286370
rect 79009 286226 79153 286370
rect 79153 286226 79212 286370
rect 78976 286176 79212 286226
rect 77081 273972 77317 274020
rect 77081 273828 77146 273972
rect 77146 273828 77290 273972
rect 77290 273828 77317 273972
rect 77081 273784 77317 273828
rect 78979 273031 79215 273072
rect 78979 272887 79016 273031
rect 79016 272887 79160 273031
rect 79160 272887 79215 273031
rect 78979 272836 79215 272887
rect 77081 260627 77317 260672
rect 77081 260483 77148 260627
rect 77148 260483 77292 260627
rect 77292 260483 77317 260627
rect 77081 260436 77317 260483
rect 78978 259680 79214 259728
rect 78978 259536 79003 259680
rect 79003 259536 79147 259680
rect 79147 259536 79214 259680
rect 78978 259492 79214 259536
rect 77080 247280 77316 247322
rect 77080 247136 77126 247280
rect 77126 247136 77270 247280
rect 77270 247136 77316 247280
rect 77080 247086 77316 247136
rect 78978 246334 79214 246374
rect 78978 246190 79017 246334
rect 79017 246190 79161 246334
rect 79161 246190 79214 246334
rect 78978 246138 79214 246190
rect 77079 233898 77315 233955
rect 77079 233754 77104 233898
rect 77104 233754 77248 233898
rect 77248 233754 77315 233898
rect 77079 233719 77315 233754
rect 78963 232952 79199 232990
rect 78963 232808 79012 232952
rect 79012 232808 79156 232952
rect 79156 232808 79199 232952
rect 78963 232754 79199 232808
rect 539228 231734 540744 233250
rect 91778 215232 92014 215254
rect 91778 215088 91818 215232
rect 91818 215088 91962 215232
rect 91962 215088 92014 215232
rect 91778 215018 92014 215088
rect 104123 215223 104359 215259
rect 104123 215079 104163 215223
rect 104163 215079 104307 215223
rect 104307 215079 104359 215223
rect 104123 215023 104359 215079
rect 117083 215101 117137 215245
rect 117137 215101 117281 215245
rect 117281 215101 117319 215245
rect 117083 215009 117319 215101
rect 129436 215183 129672 215255
rect 129436 215039 129472 215183
rect 129472 215039 129616 215183
rect 129616 215039 129672 215183
rect 129436 215019 129672 215039
rect 142741 215199 142977 215254
rect 142741 215055 142787 215199
rect 142787 215055 142931 215199
rect 142931 215055 142977 215199
rect 142741 215018 142977 215055
rect 155085 215229 155321 215256
rect 155085 215085 155127 215229
rect 155127 215085 155271 215229
rect 155271 215085 155321 215229
rect 155085 215020 155321 215085
rect 168388 215186 168624 215258
rect 168388 215042 168429 215186
rect 168429 215042 168573 215186
rect 168573 215042 168624 215186
rect 168388 215022 168624 215042
rect 180734 215217 180970 215259
rect 180734 215073 180783 215217
rect 180783 215073 180927 215217
rect 180927 215073 180970 215217
rect 180734 215023 180970 215073
rect 194025 215245 194261 215265
rect 194025 215101 194072 215245
rect 194072 215101 194216 215245
rect 194216 215101 194261 215245
rect 194025 215029 194261 215101
rect 206370 215223 206606 215258
rect 206370 215079 206430 215223
rect 206430 215079 206574 215223
rect 206574 215079 206606 215223
rect 206370 215022 206606 215079
rect 219680 215222 219916 215256
rect 219680 215078 219727 215222
rect 219727 215078 219871 215222
rect 219871 215078 219916 215222
rect 219680 215020 219916 215078
rect 232024 215113 232074 215249
rect 232074 215113 232218 215249
rect 232218 215113 232260 215249
rect 232024 215013 232260 215113
rect 245326 215241 245562 215264
rect 245326 215097 245378 215241
rect 245378 215097 245522 215241
rect 245522 215097 245562 215241
rect 245326 215028 245562 215097
rect 257668 215128 257723 215258
rect 257723 215128 257867 215258
rect 257867 215128 257904 215258
rect 257668 215022 257904 215128
rect 270987 215253 271223 215258
rect 270987 215109 271032 215253
rect 271032 215109 271176 215253
rect 271176 215109 271223 215253
rect 270987 215022 271223 215109
rect 283319 215235 283555 215261
rect 283319 215091 283375 215235
rect 283375 215091 283519 215235
rect 283519 215091 283555 215235
rect 283319 215025 283555 215091
rect 296624 215231 296860 215254
rect 296624 215087 296678 215231
rect 296678 215087 296822 215231
rect 296822 215087 296860 215231
rect 296624 215018 296860 215087
rect 308980 215238 309216 215258
rect 308980 215094 309022 215238
rect 309022 215094 309166 215238
rect 309166 215094 309216 215238
rect 308980 215022 309216 215094
rect 322257 215215 322493 215245
rect 322257 215071 322329 215215
rect 322329 215071 322473 215215
rect 322473 215071 322493 215215
rect 322257 215009 322493 215071
rect 334625 215245 334861 215256
rect 334625 215101 334673 215245
rect 334673 215101 334817 215245
rect 334817 215101 334861 215245
rect 334625 215020 334861 215101
rect 347928 215215 348164 215263
rect 347928 215071 347979 215215
rect 347979 215071 348123 215215
rect 348123 215071 348164 215215
rect 347928 215027 348164 215071
rect 360282 215227 360518 215256
rect 360282 215083 360323 215227
rect 360323 215083 360467 215227
rect 360467 215083 360518 215227
rect 360282 215020 360518 215083
rect 373576 215219 373812 215249
rect 373576 215075 373628 215219
rect 373628 215075 373772 215219
rect 373772 215075 373812 215219
rect 373576 215013 373812 215075
rect 385918 215246 386154 215259
rect 385918 215102 385973 215246
rect 385973 215102 386117 215246
rect 386117 215102 386154 215246
rect 385918 215023 386154 215102
rect 399235 215245 399471 215256
rect 399235 215101 399278 215245
rect 399278 215101 399422 215245
rect 399422 215101 399471 215245
rect 399235 215020 399471 215101
rect 411566 215211 411802 215259
rect 411566 215067 411627 215211
rect 411627 215067 411771 215211
rect 411771 215067 411802 215211
rect 411566 215023 411802 215067
rect 424885 215214 425121 215258
rect 424885 215070 424927 215214
rect 424927 215070 425071 215214
rect 425071 215070 425121 215214
rect 424885 215022 425121 215070
rect 437225 215232 437461 215258
rect 437225 215088 437275 215232
rect 437275 215088 437419 215232
rect 437419 215088 437461 215232
rect 437225 215022 437461 215088
rect 450521 215232 450757 215258
rect 450521 215088 450571 215232
rect 450571 215088 450715 215232
rect 450715 215088 450757 215232
rect 450521 215022 450757 215088
rect 462885 215219 463121 215261
rect 462885 215075 462922 215219
rect 462922 215075 463066 215219
rect 463066 215075 463121 215219
rect 462885 215025 463121 215075
rect 476187 215207 476423 215259
rect 476187 215063 476234 215207
rect 476234 215063 476378 215207
rect 476378 215063 476423 215207
rect 476187 215023 476423 215063
rect 488538 215225 488774 215259
rect 488538 215081 488575 215225
rect 488575 215081 488719 215225
rect 488719 215081 488774 215225
rect 488538 215023 488774 215081
rect 90820 213427 91056 213466
rect 90820 213283 90871 213427
rect 90871 213283 91015 213427
rect 91015 213283 91056 213427
rect 90820 213230 91056 213283
rect 103181 213425 103417 213461
rect 103181 213281 103221 213425
rect 103221 213281 103365 213425
rect 103365 213281 103417 213425
rect 103181 213225 103417 213281
rect 116145 213426 116381 213470
rect 116145 213282 116181 213426
rect 116181 213282 116325 213426
rect 116325 213282 116381 213426
rect 116145 213234 116381 213282
rect 128478 213385 128714 213458
rect 128478 213241 128524 213385
rect 128524 213241 128668 213385
rect 128668 213241 128714 213385
rect 128478 213222 128714 213241
rect 141783 213345 142019 213447
rect 141783 213211 141829 213345
rect 141829 213211 141973 213345
rect 141973 213211 142019 213345
rect 154126 213410 154362 213460
rect 154126 213266 154173 213410
rect 154173 213266 154317 213410
rect 154317 213266 154362 213410
rect 154126 213224 154362 213266
rect 167432 213371 167668 213460
rect 167432 213227 167484 213371
rect 167484 213227 167628 213371
rect 167628 213227 167668 213371
rect 167432 213224 167668 213227
rect 179791 213405 180027 213464
rect 179791 213261 179828 213405
rect 179828 213261 179972 213405
rect 179972 213261 180027 213405
rect 179791 213228 180027 213261
rect 193069 213397 193305 213464
rect 193069 213253 193138 213397
rect 193138 213253 193282 213397
rect 193282 213253 193305 213397
rect 193069 213228 193305 213253
rect 205428 213411 205664 213471
rect 205428 213267 205474 213411
rect 205474 213267 205618 213411
rect 205618 213267 205664 213411
rect 205428 213235 205664 213267
rect 218730 213412 218966 213464
rect 218730 213268 218779 213412
rect 218779 213268 218923 213412
rect 218923 213268 218966 213412
rect 218730 213228 218966 213268
rect 231074 213399 231310 213462
rect 231074 213255 231129 213399
rect 231129 213255 231273 213399
rect 231273 213255 231310 213399
rect 231074 213226 231310 213255
rect 244368 213389 244604 213458
rect 244368 213245 244428 213389
rect 244428 213245 244572 213389
rect 244572 213245 244604 213389
rect 244368 213222 244604 213245
rect 256735 213409 256971 213464
rect 256735 213265 256777 213409
rect 256777 213265 256921 213409
rect 256921 213265 256971 213409
rect 256735 213228 256971 213265
rect 270041 213390 270277 213457
rect 270041 213246 270086 213390
rect 270086 213246 270230 213390
rect 270230 213246 270277 213390
rect 270041 213221 270277 213246
rect 282367 213367 282603 213463
rect 282367 213227 282430 213367
rect 282430 213227 282574 213367
rect 282574 213227 282603 213367
rect 295678 213382 295914 213460
rect 295678 213238 295733 213382
rect 295733 213238 295877 213382
rect 295877 213238 295914 213382
rect 295678 213224 295914 213238
rect 308026 213340 308262 213453
rect 308026 213217 308081 213340
rect 308081 213217 308225 213340
rect 308225 213217 308262 213340
rect 321333 213399 321569 213458
rect 321333 213255 321379 213399
rect 321379 213255 321523 213399
rect 321523 213255 321569 213399
rect 321333 213222 321569 213255
rect 333688 213356 333924 213460
rect 333688 213224 333724 213356
rect 333724 213224 333868 213356
rect 333868 213224 333924 213356
rect 346970 213423 347206 213463
rect 346970 213279 347030 213423
rect 347030 213279 347174 213423
rect 347174 213279 347206 213423
rect 346970 213227 347206 213279
rect 359310 213411 359546 213463
rect 359310 213267 359379 213411
rect 359379 213267 359523 213411
rect 359523 213267 359546 213411
rect 359310 213227 359546 213267
rect 372639 213423 372875 213464
rect 372639 213279 372682 213423
rect 372682 213279 372826 213423
rect 372826 213279 372875 213423
rect 372639 213228 372875 213279
rect 384982 213424 385218 213464
rect 384982 213280 385029 213424
rect 385029 213280 385173 213424
rect 385173 213280 385218 213424
rect 384982 213228 385218 213280
rect 398272 213419 398508 213464
rect 398272 213275 398326 213419
rect 398326 213275 398470 213419
rect 398470 213275 398508 213419
rect 398272 213228 398508 213275
rect 410621 213419 410857 213467
rect 410621 213275 410674 213419
rect 410674 213275 410818 213419
rect 410818 213275 410857 213419
rect 410621 213231 410857 213275
rect 423941 213422 424177 213466
rect 423941 213278 423983 213422
rect 423983 213278 424127 213422
rect 424127 213278 424177 213422
rect 423941 213230 424177 213278
rect 436282 213225 436518 213461
rect 449591 213415 449827 213459
rect 449591 213271 449633 213415
rect 449633 213271 449777 213415
rect 449777 213271 449827 213415
rect 449591 213223 449827 213271
rect 461943 213413 462179 213462
rect 461943 213269 461981 213413
rect 461981 213269 462125 213413
rect 462125 213269 462179 213413
rect 461943 213226 462179 213269
rect 475223 213408 475459 213458
rect 475223 213264 475278 213408
rect 475278 213264 475422 213408
rect 475422 213264 475459 213408
rect 475223 213222 475459 213264
rect 487579 213382 487815 213463
rect 487579 213238 487626 213382
rect 487626 213238 487770 213382
rect 487770 213238 487815 213382
rect 487579 213227 487815 213238
rect 535003 213228 535239 213464
rect 569862 530707 570098 530943
rect 569603 213229 569839 213465
rect 570209 144585 570445 144821
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 8510 688382 570756 689347
rect 8510 688340 522804 688382
rect 8510 687950 512639 688340
rect 8510 687727 172302 687950
rect 8510 687491 95519 687727
rect 95755 687714 172302 687727
rect 172538 687784 512639 687950
rect 513195 687826 522804 688340
rect 523360 687826 570756 688382
rect 513195 687784 570756 687826
rect 172538 687714 570756 687784
rect 95755 687631 570756 687714
rect 95755 687625 479932 687631
rect 95755 687585 454283 687625
rect 95755 687541 223421 687585
rect 95755 687491 120844 687541
rect 8510 687305 120844 687491
rect 121080 687510 223421 687541
rect 121080 687419 216440 687510
rect 121080 687305 146501 687419
rect 8510 687183 146501 687305
rect 146737 687274 216440 687419
rect 216676 687349 223421 687510
rect 223657 687566 454283 687585
rect 223657 687540 412523 687566
rect 223657 687504 300385 687540
rect 223657 687488 274760 687504
rect 223657 687349 249091 687488
rect 216676 687274 249091 687349
rect 146737 687252 249091 687274
rect 249327 687268 274760 687488
rect 274996 687304 300385 687504
rect 300621 687505 412523 687540
rect 300621 687304 326021 687505
rect 274996 687269 326021 687304
rect 326257 687487 412523 687505
rect 326257 687269 351686 687487
rect 274996 687268 351686 687269
rect 249327 687252 351686 687268
rect 146737 687251 351686 687252
rect 351922 687449 412523 687487
rect 351922 687251 377347 687449
rect 146737 687213 377347 687251
rect 377583 687330 412523 687449
rect 412759 687556 454283 687566
rect 412759 687330 428649 687556
rect 377583 687320 428649 687330
rect 428885 687389 454283 687556
rect 454519 687395 479932 687625
rect 480168 687395 570756 687631
rect 454519 687389 570756 687395
rect 428885 687320 570756 687389
rect 377583 687213 570756 687320
rect 146737 687183 570756 687213
rect 8510 686947 570756 687183
rect 8948 530942 11348 686947
rect 8948 530706 10508 530942
rect 10744 530706 11348 530942
rect 8948 214837 11348 530706
rect 8948 214601 9916 214837
rect 10152 214601 11348 214837
rect 8948 20513 11348 214601
rect 36860 664179 541183 666579
rect 36860 542637 39260 664179
rect 36860 542401 37933 542637
rect 38169 542401 39260 542637
rect 36860 42659 39260 542401
rect 76998 434169 77398 434251
rect 76998 433933 77080 434169
rect 77316 433933 77398 434169
rect 76998 420824 77398 433933
rect 78895 433228 79295 433310
rect 78895 432992 78977 433228
rect 79213 433199 79295 433228
rect 79213 432992 79296 433199
rect 78895 432910 79296 432992
rect 76998 420588 77080 420824
rect 77316 420588 77398 420824
rect 76998 407470 77398 420588
rect 76998 407234 77080 407470
rect 77316 407234 77398 407470
rect 76998 394147 77398 407234
rect 76998 393911 77080 394147
rect 77316 393911 77398 394147
rect 76998 380781 77398 393911
rect 76998 380545 77080 380781
rect 77316 380545 77398 380781
rect 76998 367427 77398 380545
rect 76998 367191 77080 367427
rect 77316 367191 77398 367427
rect 76998 354090 77398 367191
rect 76998 353854 77080 354090
rect 77316 353854 77398 354090
rect 76998 340823 77398 353854
rect 78896 419869 79296 432910
rect 78896 419633 78978 419869
rect 79214 419633 79296 419869
rect 78896 406612 79296 419633
rect 78896 406530 79297 406612
rect 78896 406294 78979 406530
rect 79215 406294 79297 406530
rect 78896 406212 79297 406294
rect 78896 393195 79296 406212
rect 78896 392959 78978 393195
rect 79214 392959 79296 393195
rect 78896 379842 79296 392959
rect 78896 379606 78978 379842
rect 79214 379606 79296 379842
rect 78896 366568 79296 379606
rect 78896 366486 79298 366568
rect 78896 366250 78980 366486
rect 79216 366250 79298 366486
rect 78896 366168 79298 366250
rect 78896 353158 79296 366168
rect 78896 352922 78978 353158
rect 79214 352922 79296 353158
rect 76998 340741 77400 340823
rect 76998 340505 77082 340741
rect 77318 340505 77400 340741
rect 76998 340423 77400 340505
rect 76998 327458 77398 340423
rect 78896 339895 79296 352922
rect 78896 339813 79298 339895
rect 78896 339577 78980 339813
rect 79216 339577 79298 339813
rect 78896 339495 79298 339577
rect 76998 327376 77399 327458
rect 76998 327140 77081 327376
rect 77317 327140 77399 327376
rect 76998 327058 77399 327140
rect 76998 314049 77398 327058
rect 78896 326543 79296 339495
rect 78894 326461 79296 326543
rect 78894 326225 78976 326461
rect 79212 326225 79296 326461
rect 78894 326143 79296 326225
rect 76998 313813 77080 314049
rect 77316 313813 77398 314049
rect 76998 300693 77398 313813
rect 76998 300457 77080 300693
rect 77316 300457 77398 300693
rect 76998 287354 77398 300457
rect 78896 313176 79296 326143
rect 78896 313094 79297 313176
rect 78896 312858 78979 313094
rect 79215 312858 79297 313094
rect 78896 312776 79297 312858
rect 78896 299855 79296 312776
rect 78895 299773 79296 299855
rect 78895 299537 78977 299773
rect 79213 299537 79296 299773
rect 78895 299455 79296 299537
rect 76998 287118 77080 287354
rect 77316 287118 77398 287354
rect 76998 274102 77398 287118
rect 78896 286494 79296 299455
rect 78894 286412 79296 286494
rect 78894 286176 78976 286412
rect 79212 286176 79296 286412
rect 78894 286094 79296 286176
rect 76998 274020 77399 274102
rect 76998 273784 77081 274020
rect 77317 273784 77399 274020
rect 76998 273702 77399 273784
rect 76998 260754 77398 273702
rect 78896 273154 79296 286094
rect 78896 273072 79297 273154
rect 78896 272836 78979 273072
rect 79215 272836 79297 273072
rect 78896 272754 79297 272836
rect 76998 260672 77399 260754
rect 76998 260436 77081 260672
rect 77317 260436 77399 260672
rect 76998 260354 77399 260436
rect 76998 247322 77398 260354
rect 76998 247086 77080 247322
rect 77316 247086 77398 247322
rect 76998 234037 77398 247086
rect 76997 233955 77398 234037
rect 76997 233719 77079 233955
rect 77315 233719 77398 233955
rect 76997 233637 77398 233719
rect 76998 213546 77398 233637
rect 78896 259728 79296 272754
rect 78896 259492 78978 259728
rect 79214 259492 79296 259728
rect 78896 246374 79296 259492
rect 78896 246138 78978 246374
rect 79214 246138 79296 246374
rect 78896 233072 79296 246138
rect 78881 232990 79296 233072
rect 78881 232754 78963 232990
rect 79199 232754 79296 232990
rect 78881 232672 79296 232754
rect 78896 215340 79296 232672
rect 538783 233250 541183 664179
rect 538783 231734 539228 233250
rect 540744 231734 541183 233250
rect 104041 215340 104441 215341
rect 180652 215340 181052 215341
rect 193943 215340 194343 215347
rect 245244 215340 245644 215346
rect 283237 215340 283637 215343
rect 347846 215340 348246 215345
rect 385836 215340 386236 215341
rect 411484 215340 411884 215341
rect 462803 215340 463203 215343
rect 476105 215340 476505 215341
rect 488456 215340 488856 215341
rect 538783 215340 541183 231734
rect 78748 215265 541183 215340
rect 78748 215259 194025 215265
rect 78748 215254 104123 215259
rect 78748 215018 91778 215254
rect 92014 215023 104123 215254
rect 104359 215258 180734 215259
rect 104359 215256 168388 215258
rect 104359 215255 155085 215256
rect 104359 215245 129436 215255
rect 104359 215023 117083 215245
rect 92014 215018 117083 215023
rect 78748 215009 117083 215018
rect 117319 215019 129436 215245
rect 129672 215254 155085 215255
rect 129672 215019 142741 215254
rect 117319 215018 142741 215019
rect 142977 215020 155085 215254
rect 155321 215022 168388 215256
rect 168624 215023 180734 215258
rect 180970 215029 194025 215259
rect 194261 215264 541183 215265
rect 194261 215258 245326 215264
rect 194261 215029 206370 215258
rect 180970 215023 206370 215029
rect 168624 215022 206370 215023
rect 206606 215256 245326 215258
rect 206606 215022 219680 215256
rect 155321 215020 219680 215022
rect 219916 215249 245326 215256
rect 219916 215020 232024 215249
rect 142977 215018 232024 215020
rect 117319 215013 232024 215018
rect 232260 215028 245326 215249
rect 245562 215263 541183 215264
rect 245562 215261 347928 215263
rect 245562 215258 283319 215261
rect 245562 215028 257668 215258
rect 232260 215022 257668 215028
rect 257904 215022 270987 215258
rect 271223 215025 283319 215258
rect 283555 215258 347928 215261
rect 283555 215254 308980 215258
rect 283555 215025 296624 215254
rect 271223 215022 296624 215025
rect 232260 215018 296624 215022
rect 296860 215022 308980 215254
rect 309216 215256 347928 215258
rect 309216 215245 334625 215256
rect 309216 215022 322257 215245
rect 296860 215018 322257 215022
rect 232260 215013 322257 215018
rect 117319 215009 322257 215013
rect 322493 215020 334625 215245
rect 334861 215027 347928 215256
rect 348164 215261 541183 215263
rect 348164 215259 462885 215261
rect 348164 215256 385918 215259
rect 348164 215027 360282 215256
rect 334861 215020 360282 215027
rect 360518 215249 385918 215256
rect 360518 215020 373576 215249
rect 322493 215013 373576 215020
rect 373812 215023 385918 215249
rect 386154 215256 411566 215259
rect 386154 215023 399235 215256
rect 373812 215020 399235 215023
rect 399471 215023 411566 215256
rect 411802 215258 462885 215259
rect 411802 215023 424885 215258
rect 399471 215022 424885 215023
rect 425121 215022 437225 215258
rect 437461 215022 450521 215258
rect 450757 215025 462885 215258
rect 463121 215259 541183 215261
rect 463121 215025 476187 215259
rect 450757 215023 476187 215025
rect 476423 215023 488538 215259
rect 488774 215023 541183 215259
rect 450757 215022 541183 215023
rect 399471 215020 541183 215022
rect 373812 215013 541183 215020
rect 322493 215009 541183 215013
rect 78748 214940 541183 215009
rect 78896 214919 79296 214940
rect 91696 214936 92096 214940
rect 117001 214927 117401 214940
rect 129354 214937 129754 214940
rect 142659 214936 143059 214940
rect 155003 214938 155403 214940
rect 219598 214938 219998 214940
rect 231942 214931 232342 214940
rect 296542 214936 296942 214940
rect 322175 214927 322575 214940
rect 334543 214938 334943 214940
rect 360200 214938 360600 214940
rect 373494 214931 373894 214940
rect 399153 214938 399553 214940
rect 90738 213546 91138 213548
rect 116063 213546 116463 213552
rect 205346 213546 205746 213553
rect 410539 213546 410939 213549
rect 423859 213546 424259 213548
rect 76998 213471 535854 213546
rect 76998 213470 205428 213471
rect 76998 213466 116145 213470
rect 76998 213230 90820 213466
rect 91056 213461 116145 213466
rect 91056 213230 103181 213461
rect 76998 213225 103181 213230
rect 103417 213234 116145 213461
rect 116381 213464 205428 213470
rect 116381 213460 179791 213464
rect 116381 213458 154126 213460
rect 116381 213234 128478 213458
rect 103417 213225 128478 213234
rect 76998 213222 128478 213225
rect 128714 213447 154126 213458
rect 128714 213222 141783 213447
rect 76998 213211 141783 213222
rect 142019 213224 154126 213447
rect 154362 213224 167432 213460
rect 167668 213228 179791 213460
rect 180027 213228 193069 213464
rect 193305 213235 205428 213464
rect 205664 213467 535854 213471
rect 205664 213464 410621 213467
rect 205664 213235 218730 213464
rect 193305 213228 218730 213235
rect 218966 213462 256735 213464
rect 218966 213228 231074 213462
rect 167668 213226 231074 213228
rect 231310 213458 256735 213462
rect 231310 213226 244368 213458
rect 167668 213224 244368 213226
rect 142019 213222 244368 213224
rect 244604 213228 256735 213458
rect 256971 213463 372639 213464
rect 256971 213457 282367 213463
rect 256971 213228 270041 213457
rect 244604 213222 270041 213228
rect 142019 213221 270041 213222
rect 270277 213227 282367 213457
rect 282603 213460 346970 213463
rect 282603 213227 295678 213460
rect 270277 213224 295678 213227
rect 295914 213458 333688 213460
rect 295914 213453 321333 213458
rect 295914 213224 308026 213453
rect 270277 213221 308026 213224
rect 142019 213217 308026 213221
rect 308262 213222 321333 213453
rect 321569 213224 333688 213458
rect 333924 213227 346970 213460
rect 347206 213227 359310 213463
rect 359546 213228 372639 213463
rect 372875 213228 384982 213464
rect 385218 213228 398272 213464
rect 398508 213231 410621 213464
rect 410857 213466 535854 213467
rect 410857 213231 423941 213466
rect 398508 213230 423941 213231
rect 424177 213464 535854 213466
rect 424177 213463 535003 213464
rect 424177 213462 487579 213463
rect 424177 213461 461943 213462
rect 424177 213230 436282 213461
rect 398508 213228 436282 213230
rect 359546 213227 436282 213228
rect 333924 213225 436282 213227
rect 436518 213459 461943 213461
rect 436518 213225 449591 213459
rect 333924 213224 449591 213225
rect 321569 213223 449591 213224
rect 449827 213226 461943 213459
rect 462179 213458 487579 213462
rect 462179 213226 475223 213458
rect 449827 213223 475223 213226
rect 321569 213222 475223 213223
rect 475459 213227 487579 213458
rect 487815 213228 535003 213463
rect 535239 213228 535854 213464
rect 487815 213227 535854 213228
rect 475459 213222 535854 213227
rect 308262 213217 535854 213222
rect 142019 213211 535854 213217
rect 76998 213146 535854 213211
rect 103099 213143 103499 213146
rect 128396 213140 128796 213146
rect 141701 213129 142101 213146
rect 154044 213142 154444 213146
rect 167350 213142 167750 213146
rect 230992 213144 231392 213146
rect 244286 213140 244686 213146
rect 269959 213139 270359 213146
rect 282285 213145 282685 213146
rect 295596 213142 295996 213146
rect 307944 213135 308344 213146
rect 321251 213140 321651 213146
rect 333606 213142 334006 213146
rect 346888 213145 347288 213146
rect 359228 213145 359628 213146
rect 436200 213143 436600 213146
rect 449509 213141 449909 213146
rect 461861 213144 462261 213146
rect 475141 213140 475541 213146
rect 487497 213145 487897 213146
rect 538783 42659 541183 214940
rect 36860 40259 541183 42659
rect 568794 530943 571194 686947
rect 568794 530707 569862 530943
rect 570098 530707 571194 530943
rect 568794 213465 571194 530707
rect 568794 213229 569603 213465
rect 569839 213229 571194 213465
rect 568794 144821 571194 213229
rect 568794 144585 570209 144821
rect 570445 144585 571194 144821
rect 568794 20513 571194 144585
rect 8948 18113 571194 20513
use reram  reram_0
timestamp 1654740117
transform 1 0 110000 0 1 440000
box -34556 -228219 384750 119835
<< labels >>
flabel metal1 s 75892 428471 76262 428979 2 FreeSans 6108 0 0 0 V3_WL
port 1 nsew
flabel metal1 s 76076 428877 76076 428877 2 FreeSans 6108 0 0 0 V3_WL
port 1 nsew
flabel metal1 s 75878 430875 76226 431345 2 FreeSans 6108 0 0 0 V1_WL
port 2 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 4276 90 0 0 wb_clk_i
port 3 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 4276 90 0 0 wb_rst_i
port 4 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 4276 90 0 0 wbs_ack_o
port 5 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 4276 90 0 0 wbs_adr_i[0]
port 6 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 4276 90 0 0 wbs_adr_i[10]
port 7 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 4276 90 0 0 wbs_adr_i[11]
port 8 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 4276 90 0 0 wbs_adr_i[12]
port 9 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 4276 90 0 0 wbs_adr_i[13]
port 10 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 4276 90 0 0 wbs_adr_i[14]
port 11 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 4276 90 0 0 wbs_adr_i[15]
port 12 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 4276 90 0 0 wbs_adr_i[16]
port 13 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 4276 90 0 0 wbs_adr_i[17]
port 14 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 4276 90 0 0 wbs_adr_i[1]
port 15 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 4276 90 0 0 wbs_adr_i[2]
port 16 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 4276 90 0 0 wbs_adr_i[3]
port 17 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 4276 90 0 0 wbs_adr_i[4]
port 18 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 4276 90 0 0 wbs_adr_i[5]
port 19 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 4276 90 0 0 wbs_adr_i[6]
port 20 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 4276 90 0 0 wbs_adr_i[7]
port 21 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 4276 90 0 0 wbs_adr_i[8]
port 22 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 4276 90 0 0 wbs_adr_i[9]
port 23 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 4276 90 0 0 wbs_cyc_i
port 24 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 4276 90 0 0 wbs_dat_i[0]
port 25 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 4276 90 0 0 wbs_dat_i[10]
port 26 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 4276 90 0 0 wbs_dat_i[11]
port 27 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 4276 90 0 0 wbs_dat_i[12]
port 28 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 4276 90 0 0 wbs_dat_i[13]
port 29 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 4276 90 0 0 wbs_dat_i[14]
port 30 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 4276 90 0 0 wbs_dat_i[15]
port 31 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 4276 90 0 0 wbs_dat_i[16]
port 32 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 4276 90 0 0 wbs_dat_i[1]
port 33 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 4276 90 0 0 wbs_dat_i[2]
port 34 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 4276 90 0 0 wbs_dat_i[3]
port 35 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 4276 90 0 0 wbs_dat_i[4]
port 36 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 4276 90 0 0 wbs_dat_i[5]
port 37 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 4276 90 0 0 wbs_dat_i[6]
port 38 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 4276 90 0 0 wbs_dat_i[7]
port 39 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 4276 90 0 0 wbs_dat_i[8]
port 40 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 4276 90 0 0 wbs_dat_i[9]
port 41 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 4276 90 0 0 wbs_dat_o[0]
port 42 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 4276 90 0 0 wbs_dat_o[10]
port 43 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 4276 90 0 0 wbs_dat_o[11]
port 44 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 4276 90 0 0 wbs_dat_o[12]
port 45 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 4276 90 0 0 wbs_dat_o[13]
port 46 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 4276 90 0 0 wbs_dat_o[14]
port 47 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 4276 90 0 0 wbs_dat_o[15]
port 48 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 4276 90 0 0 wbs_dat_o[16]
port 49 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 4276 90 0 0 wbs_dat_o[1]
port 50 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 4276 90 0 0 wbs_dat_o[2]
port 51 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 4276 90 0 0 wbs_dat_o[3]
port 52 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 4276 90 0 0 wbs_dat_o[4]
port 53 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 4276 90 0 0 wbs_dat_o[5]
port 54 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 4276 90 0 0 wbs_dat_o[6]
port 55 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 4276 90 0 0 wbs_dat_o[7]
port 56 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 4276 90 0 0 wbs_dat_o[8]
port 57 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 4276 90 0 0 wbs_dat_o[9]
port 58 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 4276 90 0 0 wbs_sel_i[0]
port 59 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 4276 90 0 0 wbs_sel_i[1]
port 60 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 4276 90 0 0 wbs_sel_i[2]
port 61 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 4276 90 0 0 wbs_sel_i[3]
port 62 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 4276 90 0 0 wbs_stb_i
port 63 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 4276 90 0 0 wbs_we_i
port 64 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 4276 90 0 0 wbs_dat_i[17]
port 65 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 4276 90 0 0 wbs_dat_i[18]
port 66 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 4276 90 0 0 wbs_dat_i[19]
port 67 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 4276 90 0 0 wbs_adr_i[18]
port 68 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 4276 90 0 0 wbs_dat_i[20]
port 69 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 4276 90 0 0 wbs_dat_i[21]
port 70 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 4276 90 0 0 wbs_dat_i[22]
port 71 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 4276 90 0 0 wbs_dat_i[23]
port 72 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 4276 90 0 0 wbs_dat_i[24]
port 73 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 4276 90 0 0 wbs_dat_i[25]
port 74 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 4276 90 0 0 wbs_dat_i[26]
port 75 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 4276 90 0 0 wbs_dat_i[27]
port 76 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 4276 90 0 0 wbs_dat_i[28]
port 77 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 4276 90 0 0 wbs_dat_i[29]
port 78 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 4276 90 0 0 wbs_adr_i[19]
port 79 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 4276 90 0 0 wbs_dat_i[30]
port 80 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 4276 90 0 0 wbs_dat_i[31]
port 81 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 4276 90 0 0 la_oenb[0]
port 82 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 4276 90 0 0 wbs_adr_i[20]
port 83 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 4276 90 0 0 wbs_adr_i[21]
port 84 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 4276 90 0 0 wbs_adr_i[22]
port 85 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 4276 90 0 0 wbs_adr_i[23]
port 86 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 4276 90 0 0 wbs_adr_i[24]
port 87 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 4276 90 0 0 wbs_adr_i[25]
port 88 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 4276 90 0 0 wbs_adr_i[26]
port 89 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 4276 90 0 0 wbs_adr_i[27]
port 90 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 4276 90 0 0 wbs_adr_i[28]
port 91 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 4276 90 0 0 wbs_adr_i[29]
port 92 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 4276 90 0 0 la_oenb[1]
port 93 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 4276 90 0 0 wbs_adr_i[30]
port 94 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 4276 90 0 0 wbs_adr_i[31]
port 95 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 4276 90 0 0 la_oenb[2]
port 96 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 4276 90 0 0 wbs_dat_o[17]
port 97 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 4276 90 0 0 wbs_dat_o[18]
port 98 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 4276 90 0 0 wbs_dat_o[19]
port 99 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 4276 90 0 0 la_oenb[3]
port 100 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 4276 90 0 0 wbs_dat_o[20]
port 101 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 4276 90 0 0 wbs_dat_o[21]
port 102 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 4276 90 0 0 wbs_dat_o[22]
port 103 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 4276 90 0 0 wbs_dat_o[23]
port 104 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 4276 90 0 0 wbs_dat_o[24]
port 105 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 4276 90 0 0 wbs_dat_o[25]
port 106 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 4276 90 0 0 wbs_dat_o[26]
port 107 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 4276 90 0 0 wbs_dat_o[27]
port 108 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 4276 90 0 0 wbs_dat_o[28]
port 109 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 4276 90 0 0 wbs_dat_o[29]
port 110 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 4276 90 0 0 la_oenb[4]
port 111 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 4276 90 0 0 wbs_dat_o[30]
port 112 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 4276 90 0 0 wbs_dat_o[31]
port 113 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 4276 90 0 0 la_oenb[5]
port 114 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 4276 90 0 0 la_data_in[0]
port 115 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 4276 90 0 0 la_data_in[1]
port 116 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 4276 90 0 0 la_data_in[2]
port 117 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 4276 90 0 0 la_data_in[3]
port 118 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 4276 90 0 0 la_data_in[4]
port 119 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 4276 90 0 0 la_data_in[5]
port 120 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 4276 90 0 0 la_data_out[0]
port 121 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 4276 90 0 0 la_data_out[1]
port 122 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 4276 90 0 0 la_data_out[2]
port 123 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 4276 90 0 0 la_data_out[3]
port 124 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 4276 90 0 0 la_data_out[4]
port 125 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 4276 90 0 0 la_data_out[5]
port 126 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 4276 90 0 0 la_data_in[23]
port 127 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 4276 90 0 0 la_data_in[24]
port 128 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 4276 90 0 0 la_data_in[25]
port 129 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 4276 90 0 0 la_oenb[6]
port 130 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 4276 90 0 0 la_oenb[7]
port 131 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 4276 90 0 0 la_oenb[8]
port 132 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 4276 90 0 0 la_oenb[9]
port 133 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 4276 90 0 0 la_data_in[26]
port 134 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 4276 90 0 0 la_data_in[11]
port 135 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 4276 90 0 0 la_data_in[12]
port 136 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 4276 90 0 0 la_data_in[13]
port 137 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 4276 90 0 0 la_data_in[14]
port 138 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 4276 90 0 0 la_data_in[6]
port 139 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 4276 90 0 0 la_data_in[7]
port 140 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 4276 90 0 0 la_data_in[8]
port 141 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 4276 90 0 0 la_data_in[9]
port 142 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 4276 90 0 0 la_data_in[15]
port 143 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 4276 90 0 0 la_data_out[10]
port 144 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 4276 90 0 0 la_data_out[11]
port 145 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 4276 90 0 0 la_data_out[12]
port 146 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 4276 90 0 0 la_data_out[13]
port 147 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 4276 90 0 0 la_data_out[14]
port 148 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 4276 90 0 0 la_data_out[15]
port 149 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 4276 90 0 0 la_data_out[16]
port 150 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 4276 90 0 0 la_data_out[17]
port 151 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 4276 90 0 0 la_data_out[18]
port 152 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 4276 90 0 0 la_data_out[19]
port 153 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 4276 90 0 0 la_data_in[16]
port 154 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 4276 90 0 0 la_data_out[20]
port 155 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 4276 90 0 0 la_data_out[21]
port 156 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 4276 90 0 0 la_data_out[22]
port 157 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 4276 90 0 0 la_data_out[23]
port 158 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 4276 90 0 0 la_data_out[24]
port 159 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 4276 90 0 0 la_data_out[25]
port 160 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 4276 90 0 0 la_data_in[17]
port 161 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 4276 90 0 0 la_data_in[18]
port 162 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 4276 90 0 0 la_data_in[19]
port 163 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 4276 90 0 0 la_data_in[10]
port 164 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 4276 90 0 0 la_data_out[6]
port 165 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 4276 90 0 0 la_data_out[7]
port 166 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 4276 90 0 0 la_data_out[8]
port 167 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 4276 90 0 0 la_data_out[9]
port 168 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 4276 90 0 0 la_data_in[20]
port 169 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 4276 90 0 0 la_oenb[10]
port 170 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 4276 90 0 0 la_oenb[11]
port 171 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 4276 90 0 0 la_oenb[12]
port 172 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 4276 90 0 0 la_oenb[13]
port 173 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 4276 90 0 0 la_oenb[14]
port 174 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 4276 90 0 0 la_oenb[15]
port 175 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 4276 90 0 0 la_oenb[16]
port 176 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 4276 90 0 0 la_oenb[17]
port 177 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 4276 90 0 0 la_oenb[18]
port 178 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 4276 90 0 0 la_oenb[19]
port 179 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 4276 90 0 0 la_data_in[21]
port 180 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 4276 90 0 0 la_oenb[20]
port 181 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 4276 90 0 0 la_oenb[21]
port 182 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 4276 90 0 0 la_oenb[22]
port 183 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 4276 90 0 0 la_oenb[23]
port 184 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 4276 90 0 0 la_oenb[24]
port 185 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 4276 90 0 0 la_oenb[25]
port 186 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 4276 90 0 0 la_data_in[22]
port 187 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 4276 90 0 0 la_data_in[39]
port 188 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 4276 90 0 0 la_oenb[45]
port 189 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 4276 90 0 0 la_data_in[40]
port 190 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 4276 90 0 0 la_data_out[26]
port 191 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 4276 90 0 0 la_data_out[27]
port 192 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 4276 90 0 0 la_data_out[28]
port 193 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 4276 90 0 0 la_data_out[29]
port 194 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 4276 90 0 0 la_data_in[41]
port 195 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 4276 90 0 0 la_data_out[30]
port 196 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 4276 90 0 0 la_data_out[31]
port 197 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 4276 90 0 0 la_data_out[32]
port 198 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 4276 90 0 0 la_data_out[33]
port 199 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 4276 90 0 0 la_data_out[34]
port 200 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 4276 90 0 0 la_data_out[35]
port 201 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 4276 90 0 0 la_data_out[36]
port 202 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 4276 90 0 0 la_data_out[37]
port 203 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 4276 90 0 0 la_data_out[38]
port 204 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 4276 90 0 0 la_data_out[39]
port 205 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 4276 90 0 0 la_data_in[42]
port 206 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 4276 90 0 0 la_data_out[40]
port 207 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 4276 90 0 0 la_data_out[41]
port 208 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 4276 90 0 0 la_data_out[42]
port 209 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 4276 90 0 0 la_data_out[43]
port 210 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 4276 90 0 0 la_data_out[44]
port 211 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 4276 90 0 0 la_data_out[45]
port 212 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 4276 90 0 0 la_data_out[46]
port 213 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 4276 90 0 0 la_data_in[43]
port 214 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 4276 90 0 0 la_data_in[44]
port 215 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 4276 90 0 0 la_data_in[45]
port 216 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 4276 90 0 0 la_data_in[46]
port 217 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 4276 90 0 0 la_oenb[46]
port 218 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 4276 90 0 0 la_oenb[38]
port 219 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 4276 90 0 0 la_oenb[39]
port 220 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 4276 90 0 0 la_oenb[37]
port 221 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 4276 90 0 0 la_oenb[40]
port 222 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 4276 90 0 0 la_oenb[41]
port 223 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 4276 90 0 0 la_oenb[42]
port 224 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 4276 90 0 0 la_oenb[43]
port 225 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 4276 90 0 0 la_data_in[27]
port 226 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 4276 90 0 0 la_data_in[28]
port 227 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 4276 90 0 0 la_data_in[29]
port 228 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 4276 90 0 0 la_oenb[44]
port 229 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 4276 90 0 0 la_data_in[30]
port 230 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 4276 90 0 0 la_data_in[31]
port 231 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 4276 90 0 0 la_data_in[32]
port 232 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 4276 90 0 0 la_data_in[33]
port 233 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 4276 90 0 0 la_data_in[34]
port 234 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 4276 90 0 0 la_data_in[35]
port 235 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 4276 90 0 0 la_data_in[36]
port 236 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 4276 90 0 0 la_data_in[37]
port 237 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 4276 90 0 0 la_oenb[26]
port 238 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 4276 90 0 0 la_oenb[27]
port 239 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 4276 90 0 0 la_oenb[28]
port 240 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 4276 90 0 0 la_oenb[29]
port 241 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 4276 90 0 0 la_data_in[38]
port 242 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 4276 90 0 0 la_oenb[30]
port 243 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 4276 90 0 0 la_oenb[31]
port 244 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 4276 90 0 0 la_oenb[32]
port 245 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 4276 90 0 0 la_oenb[33]
port 246 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 4276 90 0 0 la_oenb[34]
port 247 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 4276 90 0 0 la_oenb[35]
port 248 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 4276 90 0 0 la_oenb[36]
port 249 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 4276 90 0 0 la_oenb[47]
port 250 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 4276 90 0 0 la_oenb[48]
port 251 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 4276 90 0 0 la_oenb[49]
port 252 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 4276 90 0 0 la_oenb[50]
port 253 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 4276 90 0 0 la_oenb[51]
port 254 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 4276 90 0 0 la_oenb[52]
port 255 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 4276 90 0 0 la_oenb[53]
port 256 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 4276 90 0 0 la_oenb[54]
port 257 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 4276 90 0 0 la_oenb[55]
port 258 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 4276 90 0 0 la_oenb[56]
port 259 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 4276 90 0 0 la_oenb[57]
port 260 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 4276 90 0 0 la_oenb[58]
port 261 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 4276 90 0 0 la_oenb[59]
port 262 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 4276 90 0 0 la_oenb[60]
port 263 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 4276 90 0 0 la_oenb[61]
port 264 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 4276 90 0 0 la_oenb[62]
port 265 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 4276 90 0 0 la_oenb[63]
port 266 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 4276 90 0 0 la_oenb[64]
port 267 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 4276 90 0 0 la_oenb[65]
port 268 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 4276 90 0 0 la_oenb[66]
port 269 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 4276 90 0 0 la_data_in[47]
port 270 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 4276 90 0 0 la_data_in[48]
port 271 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 4276 90 0 0 la_data_in[49]
port 272 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 4276 90 0 0 la_data_in[50]
port 273 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 4276 90 0 0 la_data_in[51]
port 274 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 4276 90 0 0 la_data_in[52]
port 275 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 4276 90 0 0 la_data_in[53]
port 276 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 4276 90 0 0 la_data_in[54]
port 277 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 4276 90 0 0 la_data_in[55]
port 278 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 4276 90 0 0 la_data_in[56]
port 279 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 4276 90 0 0 la_data_in[57]
port 280 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 4276 90 0 0 la_data_in[58]
port 281 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 4276 90 0 0 la_data_in[59]
port 282 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 4276 90 0 0 la_data_in[60]
port 283 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 4276 90 0 0 la_data_in[61]
port 284 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 4276 90 0 0 la_data_in[62]
port 285 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 4276 90 0 0 la_data_in[63]
port 286 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 4276 90 0 0 la_data_out[47]
port 287 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 4276 90 0 0 la_data_out[48]
port 288 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 4276 90 0 0 la_data_out[49]
port 289 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 4276 90 0 0 la_data_in[64]
port 290 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 4276 90 0 0 la_data_out[50]
port 291 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 4276 90 0 0 la_data_out[51]
port 292 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 4276 90 0 0 la_data_out[52]
port 293 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 4276 90 0 0 la_data_out[53]
port 294 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 4276 90 0 0 la_data_out[54]
port 295 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 4276 90 0 0 la_data_out[55]
port 296 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 4276 90 0 0 la_data_out[56]
port 297 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 4276 90 0 0 la_data_out[57]
port 298 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 4276 90 0 0 la_data_out[58]
port 299 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 4276 90 0 0 la_data_out[59]
port 300 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 4276 90 0 0 la_data_in[65]
port 301 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 4276 90 0 0 la_data_out[60]
port 302 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 4276 90 0 0 la_data_out[61]
port 303 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 4276 90 0 0 la_data_out[62]
port 304 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 4276 90 0 0 la_data_out[63]
port 305 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 4276 90 0 0 la_data_out[64]
port 306 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 4276 90 0 0 la_data_out[65]
port 307 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 4276 90 0 0 la_data_out[66]
port 308 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 4276 90 0 0 la_data_out[67]
port 309 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 4276 90 0 0 la_data_in[66]
port 310 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 4276 90 0 0 la_data_in[67]
port 311 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 4276 90 0 0 la_data_in[72]
port 312 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 4276 90 0 0 la_data_in[73]
port 313 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 4276 90 0 0 la_data_in[74]
port 314 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 4276 90 0 0 la_data_in[75]
port 315 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 4276 90 0 0 la_data_in[76]
port 316 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 4276 90 0 0 la_data_in[77]
port 317 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 4276 90 0 0 la_data_in[78]
port 318 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 4276 90 0 0 la_data_in[79]
port 319 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 4276 90 0 0 la_data_in[80]
port 320 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 4276 90 0 0 la_data_in[81]
port 321 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 4276 90 0 0 la_data_in[82]
port 322 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 4276 90 0 0 la_data_in[83]
port 323 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 4276 90 0 0 la_data_in[84]
port 324 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 4276 90 0 0 la_data_in[85]
port 325 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 4276 90 0 0 la_data_in[86]
port 326 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 4276 90 0 0 la_data_in[87]
port 327 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 4276 90 0 0 la_data_in[69]
port 328 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 4276 90 0 0 la_oenb[67]
port 329 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 4276 90 0 0 la_oenb[68]
port 330 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 4276 90 0 0 la_oenb[69]
port 331 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 4276 90 0 0 la_oenb[70]
port 332 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 4276 90 0 0 la_oenb[71]
port 333 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 4276 90 0 0 la_oenb[72]
port 334 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 4276 90 0 0 la_oenb[73]
port 335 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 4276 90 0 0 la_oenb[74]
port 336 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 4276 90 0 0 la_oenb[75]
port 337 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 4276 90 0 0 la_oenb[76]
port 338 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 4276 90 0 0 la_oenb[77]
port 339 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 4276 90 0 0 la_oenb[78]
port 340 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 4276 90 0 0 la_oenb[79]
port 341 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 4276 90 0 0 la_oenb[80]
port 342 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 4276 90 0 0 la_oenb[81]
port 343 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 4276 90 0 0 la_oenb[82]
port 344 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 4276 90 0 0 la_oenb[83]
port 345 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 4276 90 0 0 la_oenb[84]
port 346 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 4276 90 0 0 la_oenb[85]
port 347 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 4276 90 0 0 la_oenb[86]
port 348 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 4276 90 0 0 la_oenb[87]
port 349 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 4276 90 0 0 la_data_out[68]
port 350 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 4276 90 0 0 la_data_out[69]
port 351 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 4276 90 0 0 la_data_in[70]
port 352 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 4276 90 0 0 la_data_out[70]
port 353 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 4276 90 0 0 la_data_out[71]
port 354 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 4276 90 0 0 la_data_out[72]
port 355 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 4276 90 0 0 la_data_out[73]
port 356 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 4276 90 0 0 la_data_out[74]
port 357 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 4276 90 0 0 la_data_out[75]
port 358 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 4276 90 0 0 la_data_out[76]
port 359 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 4276 90 0 0 la_data_out[77]
port 360 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 4276 90 0 0 la_data_out[78]
port 361 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 4276 90 0 0 la_data_out[79]
port 362 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 4276 90 0 0 la_data_in[71]
port 363 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 4276 90 0 0 la_data_out[80]
port 364 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 4276 90 0 0 la_data_out[81]
port 365 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 4276 90 0 0 la_data_out[82]
port 366 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 4276 90 0 0 la_data_out[83]
port 367 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 4276 90 0 0 la_data_out[84]
port 368 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 4276 90 0 0 la_data_out[85]
port 369 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 4276 90 0 0 la_data_out[86]
port 370 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 4276 90 0 0 la_data_out[87]
port 371 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 4276 90 0 0 la_data_in[68]
port 372 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 4276 90 0 0 la_oenb[88]
port 373 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 4276 90 0 0 la_oenb[89]
port 374 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 4276 90 0 0 la_oenb[90]
port 375 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 4276 90 0 0 la_oenb[91]
port 376 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 4276 90 0 0 la_oenb[92]
port 377 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 4276 90 0 0 la_oenb[93]
port 378 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 4276 90 0 0 la_oenb[94]
port 379 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 4276 90 0 0 la_oenb[95]
port 380 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 4276 90 0 0 la_oenb[96]
port 381 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 4276 90 0 0 la_oenb[97]
port 382 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 4276 90 0 0 la_oenb[98]
port 383 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 4276 90 0 0 la_oenb[99]
port 384 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 4276 90 0 0 la_data_in[101]
port 385 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 4276 90 0 0 la_data_in[102]
port 386 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 4276 90 0 0 la_data_in[103]
port 387 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 4276 90 0 0 la_data_in[104]
port 388 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 4276 90 0 0 la_data_in[105]
port 389 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 4276 90 0 0 la_data_in[106]
port 390 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 4276 90 0 0 la_data_in[107]
port 391 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 4276 90 0 0 la_data_in[108]
port 392 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 4276 90 0 0 la_data_in[100]
port 393 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 4276 90 0 0 la_data_in[90]
port 394 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 4276 90 0 0 la_data_in[91]
port 395 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 4276 90 0 0 la_data_in[92]
port 396 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 4276 90 0 0 la_data_in[93]
port 397 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 4276 90 0 0 la_data_in[94]
port 398 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 4276 90 0 0 la_data_in[95]
port 399 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 4276 90 0 0 la_data_in[96]
port 400 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 4276 90 0 0 la_data_in[97]
port 401 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 4276 90 0 0 la_data_in[98]
port 402 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 4276 90 0 0 la_data_in[99]
port 403 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 4276 90 0 0 la_data_out[100]
port 404 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 4276 90 0 0 la_data_out[101]
port 405 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 4276 90 0 0 la_data_out[102]
port 406 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 4276 90 0 0 la_data_out[103]
port 407 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 4276 90 0 0 la_data_out[104]
port 408 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 4276 90 0 0 la_data_out[105]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 4276 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 4276 90 0 0 la_data_out[106]
port 411 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 4276 90 0 0 la_data_out[94]
port 412 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 4276 90 0 0 la_data_out[107]
port 413 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 4276 90 0 0 la_data_out[95]
port 414 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 4276 90 0 0 la_data_out[96]
port 415 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 4276 90 0 0 la_data_out[108]
port 416 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 4276 90 0 0 la_data_out[97]
port 417 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 4276 90 0 0 la_data_out[98]
port 418 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 4276 90 0 0 la_data_out[99]
port 419 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 4276 90 0 0 la_data_out[92]
port 420 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 4276 90 0 0 la_oenb[100]
port 421 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 4276 90 0 0 la_oenb[101]
port 422 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 4276 90 0 0 la_oenb[102]
port 423 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 4276 90 0 0 la_oenb[103]
port 424 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 4276 90 0 0 la_oenb[104]
port 425 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 4276 90 0 0 la_oenb[105]
port 426 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 4276 90 0 0 la_oenb[106]
port 427 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 4276 90 0 0 la_oenb[107]
port 428 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 4276 90 0 0 la_data_in[88]
port 429 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 4276 90 0 0 la_data_in[89]
port 430 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 4276 90 0 0 la_data_out[88]
port 431 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 4276 90 0 0 la_data_out[89]
port 432 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 4276 90 0 0 la_data_out[90]
port 433 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 4276 90 0 0 la_data_out[91]
port 434 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 4276 90 0 0 la_data_in[119]
port 435 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 4276 90 0 0 la_data_out[120]
port 436 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 4276 90 0 0 la_data_out[121]
port 437 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 4276 90 0 0 la_data_out[122]
port 438 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 4276 90 0 0 la_data_in[116]
port 439 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 4276 90 0 0 la_data_in[117]
port 440 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 4276 90 0 0 la_data_out[123]
port 441 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 4276 90 0 0 la_data_in[112]
port 442 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 4276 90 0 0 la_data_out[124]
port 443 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 4276 90 0 0 la_data_out[125]
port 444 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 4276 90 0 0 la_data_out[126]
port 445 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 4276 90 0 0 la_data_out[127]
port 446 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 4276 90 0 0 la_data_in[118]
port 447 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 4276 90 0 0 la_oenb[109]
port 448 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 4276 90 0 0 la_data_in[120]
port 449 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 4276 90 0 0 la_oenb[110]
port 450 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 4276 90 0 0 la_data_in[121]
port 451 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 4276 90 0 0 la_oenb[111]
port 452 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 4276 90 0 0 la_oenb[112]
port 453 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 4276 90 0 0 la_oenb[113]
port 454 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 4276 90 0 0 la_oenb[114]
port 455 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 4276 90 0 0 la_oenb[115]
port 456 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 4276 90 0 0 la_oenb[116]
port 457 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 4276 90 0 0 la_oenb[117]
port 458 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 4276 90 0 0 la_oenb[118]
port 459 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 4276 90 0 0 la_oenb[119]
port 460 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 4276 90 0 0 la_data_in[122]
port 461 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 4276 90 0 0 la_data_in[123]
port 462 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 4276 90 0 0 la_oenb[120]
port 463 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 4276 90 0 0 la_oenb[121]
port 464 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 4276 90 0 0 la_oenb[122]
port 465 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 4276 90 0 0 la_oenb[123]
port 466 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 4276 90 0 0 la_oenb[124]
port 467 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 4276 90 0 0 la_oenb[125]
port 468 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 4276 90 0 0 la_oenb[126]
port 469 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 4276 90 0 0 la_oenb[127]
port 470 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 4276 90 0 0 la_data_in[124]
port 471 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 4276 90 0 0 la_data_in[125]
port 472 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 4276 90 0 0 la_data_in[126]
port 473 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 4276 90 0 0 la_data_in[127]
port 474 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 4276 90 0 0 la_data_out[110]
port 475 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 4276 90 0 0 user_clock2
port 476 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 4276 90 0 0 user_irq[0]
port 477 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 4276 90 0 0 la_data_in[113]
port 478 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 4276 90 0 0 user_irq[1]
port 479 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 4276 90 0 0 la_data_in[114]
port 480 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 4276 90 0 0 user_irq[2]
port 481 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 4276 90 0 0 la_data_out[111]
port 482 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 4276 90 0 0 la_data_out[112]
port 483 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 4276 90 0 0 la_data_out[109]
port 484 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 4276 90 0 0 la_data_in[109]
port 485 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 4276 90 0 0 la_data_out[113]
port 486 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 4276 90 0 0 la_data_in[110]
port 487 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 4276 90 0 0 la_data_out[114]
port 488 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 4276 90 0 0 la_oenb[108]
port 489 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 4276 90 0 0 la_data_out[115]
port 490 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 4276 90 0 0 la_data_out[116]
port 491 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 4276 90 0 0 la_data_in[111]
port 492 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 4276 90 0 0 la_data_out[117]
port 493 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 4276 90 0 0 la_data_in[115]
port 494 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 4276 90 0 0 la_data_out[118]
port 495 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 4276 90 0 0 la_data_out[119]
port 496 nsew
flabel mvpsubdiff s 76026 431246 76026 431246 2 FreeSans 6108 0 0 0 V1_WL
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 7326 180 0 0 io_analog[4]
port 497 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 7326 180 0 0 io_analog[4]
port 497 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 7326 180 0 0 io_analog[5]
port 498 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 7326 180 0 0 io_analog[5]
port 498 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 7326 180 0 0 io_analog[6]
port 499 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 7326 180 0 0 io_analog[6]
port 499 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 7326 180 0 0 io_analog[4]
port 497 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 7326 180 0 0 io_analog[4]
port 497 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 4276 0 0 0 gpio_analog[2]
port 500 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 4276 0 0 0 gpio_analog[3]
port 501 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 4276 0 0 0 gpio_analog[4]
port 502 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 4276 0 0 0 gpio_analog[5]
port 503 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 4276 0 0 0 gpio_analog[6]
port 504 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 4276 0 0 0 gpio_noesd[2]
port 505 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 4276 0 0 0 gpio_noesd[3]
port 506 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 4276 0 0 0 gpio_noesd[4]
port 507 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 4276 0 0 0 gpio_noesd[5]
port 508 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 4276 0 0 0 gpio_noesd[6]
port 509 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 4276 0 0 0 io_analog[0]
port 510 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 7326 180 0 0 io_analog[1]
port 511 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 7326 180 0 0 io_analog[2]
port 512 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 7326 180 0 0 io_analog[3]
port 513 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 7326 180 0 0 io_clamp_high[0]
port 514 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 7326 180 0 0 io_clamp_low[0]
port 515 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 4276 0 0 0 io_in[10]
port 516 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 4276 0 0 0 io_in[11]
port 517 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 4276 0 0 0 io_in[12]
port 518 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 4276 0 0 0 io_in[13]
port 519 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 4276 0 0 0 io_in[9]
port 520 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 4276 0 0 0 io_in_3v3[10]
port 521 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 4276 0 0 0 io_in_3v3[11]
port 522 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 4276 0 0 0 io_in_3v3[12]
port 523 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 4276 0 0 0 io_in_3v3[13]
port 524 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 4276 0 0 0 io_in_3v3[9]
port 525 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 4276 0 0 0 io_oeb[10]
port 526 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 4276 0 0 0 io_oeb[11]
port 527 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 4276 0 0 0 io_oeb[12]
port 528 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 4276 0 0 0 io_oeb[13]
port 529 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 4276 0 0 0 io_oeb[9]
port 530 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 4276 0 0 0 io_out[10]
port 531 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 4276 0 0 0 io_out[11]
port 532 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 4276 0 0 0 io_out[12]
port 533 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 4276 0 0 0 io_out[13]
port 534 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 4276 0 0 0 io_out[9]
port 535 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 4276 0 0 0 vccd1
port 536 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 4276 0 0 0 vccd1
port 536 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 4276 0 0 0 vdda1
port 537 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 4276 0 0 0 vdda1
port 537 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 7326 180 0 0 vssa1
port 538 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 7326 180 0 0 vssa1
port 538 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 7326 180 0 0 io_analog[6]
port 499 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 7326 180 0 0 io_analog[6]
port 499 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 7326 180 0 0 io_analog[5]
port 498 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 7326 180 0 0 io_analog[5]
port 498 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 4276 0 0 0 io_in[16]
port 539 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 4276 0 0 0 io_in[17]
port 540 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 4276 0 0 0 gpio_analog[9]
port 541 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 4276 0 0 0 gpio_noesd[10]
port 542 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 7326 180 0 0 io_analog[7]
port 543 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 4276 0 0 0 io_in_3v3[14]
port 544 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 4276 0 0 0 io_in_3v3[15]
port 545 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 4276 0 0 0 io_in_3v3[16]
port 546 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 4276 0 0 0 io_in_3v3[17]
port 547 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 7326 180 0 0 io_analog[8]
port 548 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 7326 180 0 0 io_analog[9]
port 549 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 4276 0 0 0 gpio_noesd[7]
port 550 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 4276 0 0 0 io_oeb[14]
port 551 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 4276 0 0 0 io_oeb[15]
port 552 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 4276 0 0 0 io_oeb[16]
port 553 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 4276 0 0 0 io_oeb[17]
port 554 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 4276 0 0 0 gpio_noesd[8]
port 555 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 7326 180 0 0 io_clamp_high[1]
port 556 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 7326 180 0 0 io_clamp_high[2]
port 557 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 4276 0 0 0 gpio_noesd[9]
port 558 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 7326 180 0 0 io_clamp_low[1]
port 559 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 4276 0 0 0 io_out[14]
port 560 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 4276 0 0 0 io_out[15]
port 561 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 4276 0 0 0 io_out[16]
port 562 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 4276 0 0 0 io_out[17]
port 563 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 7326 180 0 0 io_clamp_low[2]
port 564 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 4276 0 0 0 gpio_analog[10]
port 565 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 4276 0 0 0 io_analog[10]
port 566 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 4276 0 0 0 vccd2
port 567 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 4276 0 0 0 vccd2
port 567 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 4276 0 0 0 gpio_analog[7]
port 568 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 4276 0 0 0 gpio_analog[8]
port 569 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 4276 0 0 0 io_in[14]
port 570 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 4276 0 0 0 io_in[15]
port 571 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 4276 0 0 0 vssa2
port 572 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 4276 0 0 0 vssa2
port 572 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 4276 0 0 0 io_in_3v3[24]
port 573 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 4276 0 0 0 io_in_3v3[25]
port 574 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 4276 0 0 0 io_in_3v3[26]
port 575 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 4276 0 0 0 gpio_analog[16]
port 576 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 4276 0 0 0 gpio_analog[17]
port 577 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 4276 0 0 0 gpio_analog[11]
port 578 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 4276 0 0 0 gpio_analog[12]
port 579 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 4276 0 0 0 gpio_noesd[11]
port 580 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 4276 0 0 0 io_in[18]
port 581 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 4276 0 0 0 io_in[19]
port 582 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 4276 0 0 0 io_in[20]
port 583 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 4276 0 0 0 io_in[21]
port 584 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 4276 0 0 0 io_oeb[18]
port 585 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 4276 0 0 0 io_oeb[19]
port 586 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 4276 0 0 0 io_oeb[20]
port 587 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 4276 0 0 0 io_oeb[21]
port 588 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 4276 0 0 0 io_oeb[22]
port 589 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 4276 0 0 0 io_oeb[23]
port 590 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 4276 0 0 0 io_oeb[24]
port 591 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 4276 0 0 0 io_oeb[25]
port 592 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 4276 0 0 0 io_oeb[26]
port 593 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 4276 0 0 0 io_in[22]
port 594 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 4276 0 0 0 io_in[23]
port 595 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 4276 0 0 0 io_in[24]
port 596 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 4276 0 0 0 io_in[25]
port 597 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 4276 0 0 0 io_in[26]
port 598 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 4276 0 0 0 gpio_noesd[12]
port 599 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 4276 0 0 0 gpio_noesd[13]
port 600 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 4276 0 0 0 gpio_noesd[14]
port 601 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 4276 0 0 0 gpio_noesd[15]
port 602 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 4276 0 0 0 io_out[18]
port 603 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 4276 0 0 0 io_out[19]
port 604 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 4276 0 0 0 io_out[20]
port 605 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 4276 0 0 0 io_out[21]
port 606 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 4276 0 0 0 io_out[22]
port 607 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 4276 0 0 0 io_out[23]
port 608 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 4276 0 0 0 io_out[24]
port 609 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 4276 0 0 0 io_out[25]
port 610 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 4276 0 0 0 io_out[26]
port 611 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 4276 0 0 0 gpio_noesd[16]
port 612 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 4276 0 0 0 gpio_noesd[17]
port 613 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 4276 0 0 0 gpio_analog[13]
port 614 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 4276 0 0 0 gpio_analog[14]
port 615 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 4276 0 0 0 gpio_analog[15]
port 616 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 4276 0 0 0 io_in_3v3[18]
port 617 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 4276 0 0 0 io_in_3v3[19]
port 618 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 4276 0 0 0 vdda2
port 619 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 4276 0 0 0 vdda2
port 619 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 4276 0 0 0 io_in_3v3[20]
port 620 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 4276 0 0 0 io_in_3v3[21]
port 621 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 4276 0 0 0 io_in_3v3[22]
port 622 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 4276 0 0 0 io_in_3v3[23]
port 623 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 4276 0 0 0 vssd2
port 624 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 4276 0 0 0 vssd2
port 624 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 4276 0 0 0 vssa1
port 538 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 4276 0 0 0 vssa1
port 538 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 4276 0 0 0 vdda1
port 537 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 4276 0 0 0 vdda1
port 537 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 4276 0 0 0 io_in_3v3[6]
port 625 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 4276 0 0 0 io_in_3v3[7]
port 626 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 4276 0 0 0 io_in_3v3[8]
port 627 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 4276 0 0 0 io_in[1]
port 628 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 4276 0 0 0 io_oeb[0]
port 629 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 4276 0 0 0 gpio_noesd[0]
port 630 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 4276 0 0 0 io_in[2]
port 631 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 4276 0 0 0 io_in[3]
port 632 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 4276 0 0 0 io_in[4]
port 633 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 4276 0 0 0 io_in[5]
port 634 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 4276 0 0 0 io_out[1]
port 635 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 4276 0 0 0 io_in[6]
port 636 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 4276 0 0 0 io_in_3v3[1]
port 637 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 4276 0 0 0 io_in[7]
port 638 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 4276 0 0 0 io_in[8]
port 639 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 4276 0 0 0 gpio_analog[0]
port 640 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 4276 0 0 0 io_oeb[1]
port 641 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 4276 0 0 0 io_in_3v3[0]
port 642 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 4276 0 0 0 io_out[2]
port 643 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 4276 0 0 0 io_out[3]
port 644 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 4276 0 0 0 io_out[4]
port 645 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 4276 0 0 0 io_out[5]
port 646 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 4276 0 0 0 io_out[6]
port 647 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 4276 0 0 0 io_out[7]
port 648 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 4276 0 0 0 io_out[8]
port 649 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 4276 0 0 0 gpio_analog[1]
port 650 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 4276 0 0 0 gpio_noesd[1]
port 651 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 4276 0 0 0 io_in[0]
port 652 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 4276 0 0 0 io_in_3v3[2]
port 653 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 4276 0 0 0 io_in_3v3[3]
port 654 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 4276 0 0 0 io_in_3v3[4]
port 655 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 4276 0 0 0 io_oeb[2]
port 656 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 4276 0 0 0 io_oeb[3]
port 657 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 4276 0 0 0 io_oeb[4]
port 658 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 4276 0 0 0 io_oeb[5]
port 659 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 4276 0 0 0 io_oeb[6]
port 660 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 4276 0 0 0 io_oeb[7]
port 661 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 4276 0 0 0 io_oeb[8]
port 662 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 4276 0 0 0 vssd1
port 663 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 4276 0 0 0 vssd1
port 663 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 4276 0 0 0 io_in_3v3[5]
port 664 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 4276 0 0 0 io_out[0]
port 665 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 7326 180 0 0 io_analog[4]
port 497 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 7326 180 0 0 io_analog[4]
port 497 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 7326 180 0 0 io_analog[5]
port 498 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 7326 180 0 0 io_analog[5]
port 498 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 7326 180 0 0 io_analog[6]
port 499 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 7326 180 0 0 io_analog[6]
port 499 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
